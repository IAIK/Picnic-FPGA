library ieee;
use ieee.std_logic_1164.all;

library work;

package lowmc_pkg is
  constant N : integer := 128;
  constant K : integer := 128;
  constant M : integer := 10;
  constant R : integer := 20;
  constant S : integer := 30;

  type T_NK_MATRIX is array(0 to N - 1) of std_logic_vector(K - 1 downto 0);
  type T_NN_MATRIX is array(0 to N - 1) of std_logic_vector(N - 1 downto 0);
  type T_SK_MATRIX is array(0 to S - 1) of std_logic_vector(K - 1 downto 0);
  type T_SN_MATRIX is array(0 to S - 1) of std_logic_vector(N - 1 downto 0);
  type T_NSS_MATRIX is array(0 to (N - S) - 1) of std_logic_vector(S - 1 downto 0);
  type T_RS_MATRIX is array(0 to R - 1) of std_logic_vector(S - 1 downto 0);

  type T_KMATRIX is array (0 to R - 1) of T_SK_MATRIX;
  type T_ZMATRIX is array (0 to R - 2) of T_SN_MATRIX;
  type T_RMATRIX is array (0 to R - 2) of T_NSS_MATRIX;

  constant K0 : T_NK_MATRIX := (
      x"fb126337ed0ffbf2e4389aac9149432e",
      x"a216877dc9614af485edaa32f8f9fc28",
      x"67b0aec751ded3c7fed3b03634447822",
      x"1ffe172d815e9eff9449c29f8d9100a3",
      x"124cbc5eb7bb30248d95333a7e9014ab",
      x"ab8df29ec3528a45f515863b4b6cebd8",
      x"67aa2a15203866be7740574fbe22c4d8",
      x"0012c7b7d61b5993bed9d6476a0465a8",
      x"4547ea59e55c31b5686326707301fda5",
      x"1921b4c7fcd32cd2f302693fcb3ab4c9",
      x"13283c51db8b4bb7667db6e8f922a7bc",
      x"940d6cae905019d5153814bfa1f8b488",
      x"cae62c1a9434247e2ab99722ee59c8be",
      x"df7226935c6d09fd1de9e3922b268a58",
      x"6c16fd1887db4f0e11ceaecabaaaf5cb",
      x"c79611ee55a26e6c005815f825d49b3c",
      x"43498ed8f5c297e0502d5a406a1e6c50",
      x"cc583650117553374874594e66db175c",
      x"aa44dcdab477cb6769591483ae9438db",
      x"a44ecf9fe772f5eb663e256d64dc07c7",
      x"91dfc7e9651fdd64f9ba26632bd7dbd5",
      x"2d25b07947adfe4c10845f4650acbcb1",
      x"f908ca1ee240144e99c8ed66fd1b1316",
      x"9a103eca8cc6143c6677b79ed93eefad",
      x"d0226093e30063a930561820af6370c8",
      x"d112abfde53efb6fdc7032ed10c8ce11",
      x"d1caa04dacd7ab1f65e90851e18a3606",
      x"797f81a6308d057450c5d9b1029e425f",
      x"c4174e16e1c3af85c13fe8315df66c71",
      x"dab2eb8443a0e0a169eba6668472019a",
      x"f1a547aefb8b17b5077be24d1fab367f",
      x"7a913da94dc25dd6ae5a1fb1c0382345",
      x"3a3b1e7b0e91f8b1b874ea6fcc0bddf6",
      x"a16f6d344ea82e581c9f5862f65160cf",
      x"9b564bbece1cdb8da0b366a6d36b5c24",
      x"ac92cef46f6359607f138f7d9260372f",
      x"c36935b703ada0f862eea1cb0bd36b7b",
      x"1b3500c999b03dd3f2eccefd9bea35db",
      x"7333599d72ef122b108b52d58288239f",
      x"8848c586c7ee526d885fd16d3ae55954",
      x"77c2cf5adcfcd8e261f2add2aa4674a5",
      x"4b4e746a6cd6b5b0e06c89adfa004203",
      x"d8a73df034c0b2a5ae54a95ab0cfd34e",
      x"7129f8a73213b022fd0d02b470d59a11",
      x"b6aa121739c7e845eadc3db63ed29daf",
      x"fb63b0c719e8e3561874b9bc7d43b785",
      x"e61854153f346f9a13942cef20d2723b",
      x"155bcac97153967f00115048603bf1ae",
      x"877cb6a8e89ca3cddd2a562de758a5dc",
      x"185968989c1d86b25cad3c34a59b5419",
      x"af1dbdb80f5daed18cb1f2da9a99d8c7",
      x"dac33739271995e92180253961730f17",
      x"18a78da5cfe4b173e61c884b6980c77e",
      x"1facfc3609902cfe25bef826fb636b6b",
      x"6a744c36d26f6798ded507b05a770881",
      x"869ecce165d6f507fdc2efc40a9a6df8",
      x"99621ab0a3470976b2eead2b9fd83e81",
      x"4b6451eb6d67b9a3fcef89a225d68563",
      x"148dd7fbdc1ec30a87e037fb0b5f8c0d",
      x"ddf0e8d97acf8052b28129e275324db7",
      x"a12ee70f29635f1ce3857157feb9ddff",
      x"42498baa4706420d03daaab9ddd1716b",
      x"6d5233d6e214c6cd86fe99a70e617e9d",
      x"d80dec33028dc58a1a5b70acc767e8c8",
      x"c49f9ee9258e6d10bc6e371879e33f52",
      x"f17a25f6b784cc1df80e5c5c45adf907",
      x"d7774eeeb2023df7b53e265ce3e7df69",
      x"ab24cde1d3efc82d4f522d7dd904e6bc",
      x"a9ac5f83e320bc129bef20f9834506aa",
      x"d9586b72bd7a6e11e9c1c5c05c35377c",
      x"76113a1e7eb738c6abb4b38f8f35d628",
      x"f1152f66ad2d4d6893b66b89b7f036e7",
      x"c34e163b5df24aa9f77ca933428d6b87",
      x"1f227604ed461186e5349b31010a3a81",
      x"eaf3f81da6390e624975e396809984cd",
      x"0baed6fe121d178e155b6bc5e0530e04",
      x"b094ba94380726a06fe1569cc15037b0",
      x"3272f43bd5a707e262d9a8607d326836",
      x"74c4b0a12413604f70c65911eacd9bea",
      x"e07204bdd0d4a156adea009f6c6c1bf9",
      x"a94e4c665ba16e6477dc3402011d5624",
      x"e2842ac82c32c258993344326950914e",
      x"4e95767b787bd7edac11da37431eeaeb",
      x"875ee0dbaaa5a2c086e02dc09d40bda0",
      x"528f15f12fbc6151782309ab7799d35a",
      x"3fa1b6bd90bd41c2557627ab1a51425b",
      x"9463c9b69af14fb9c8ee7de0df78239c",
      x"1f0948278fb4b545ff87b4ecf3bd4d28",
      x"3cd8722b811524cf218a68447a40046f",
      x"c53d438812d2505713c3e6bf0bedae3f",
      x"5f417dae0d24c42eac7fdf162a3dc30c",
      x"59eb2b0c35894dc8af82412ffc39cae8",
      x"136043192d7b535bc180fbe50179ee3d",
      x"bee3c3c0f8a1929315c4718e5f11a4ad",
      x"e9f65681d1f4df1900da0f0bbd896b5e",
      x"30f583463ac6e1b57fd8c961d82591d9",
      x"48117d039afcbc2f8f8d20384f20bb24",
      x"3ee2494529841deba51f588fe58afeda",
      x"4e24162730965863d383e751489c358b",
      x"a922c1b6abfde633d8b4972364632e7c",
      x"ea4bbb24664639c8f69c2ad82c2942d4",
      x"3a18d07f2583d80ec0a7d9505f059aac",
      x"014d0eae53b7deb42987d554ff9dcc96",
      x"5b022239191054a5f9bf0dd0ea492015",
      x"726f052c760684fc5f8685ecdbc9cd99",
      x"75a77542d236a0a9987a180734610aa4",
      x"6899842c62755634080bc87bdd498a14",
      x"d93abb98c1a05eb027549b6906fef167",
      x"f1b5230ecac6986a02183f931202b470",
      x"a6eef93fcea9abff424faba6f73d2582",
      x"fd0e1037f88c0599a74f7e986bbe21d8",
      x"8c5be1f28d86ebf70c44e62e11b645a9",
      x"244e2834c29c1c87ed012530b302f7af",
      x"c347ae2058341fe84f76b117aa42dc8e",
      x"7363bbc6d29ae3eb58ce76d3f1f1813a",
      x"503ecbc90405f13a84c34620c4081ad8",
      x"4931fb6a84b25f8afb56d1515e3002b6",
      x"4d95b94014e1127a4c011fe406382446",
      x"a8c156ea081feec035d3650fbf454a18",
      x"658715c518fd0cd544d121e1c4f1f38d",
      x"3c2b1683311a804128c22273d9ba3a82",
      x"bc51ce30cab9ab8ebbfba740546efaff",
      x"910fb2b3cdd0ff0746a01e1ac630ae49",
      x"ad771374a75d78344ccd812b1601e0a6",
      x"501bb443ae45feb672f3dc4d68ceaad5",
      x"a3563023f7868463ed42a4feaf6ce75f",
      x"218c997316b9c3c5e6da4ff0f21320d9",
      x"6ba789fdfdb5e524b0b76898156f090e"
  );

  constant KMATRIX : T_KMATRIX := (
    (
      x"d69a7d0500f0be1a0afa96e582f026dd",
      x"ae0a095093afe4ed95996a75b86eb0c9",
      x"0f8531f7e9241696fd6310ea5d69543c",
      x"efa75ed4a280b683fd71c13b6661bf2c",
      x"95e965a594363622d7373e12850aa9ae",
      x"2c5e1b0fa9bd45cde1230e5bd304da0c",
      x"6afb80843997b9084b6dbdceccb1b9b9",
      x"f36aa16e2dea00e2a890e7613822e79f",
      x"32e601749fa50ebec137310dbe514ca5",
      x"778cd8353d2242ee038dd5177b470ee1",
      x"60510da3f88fa88ff6329db8e6aaaf16",
      x"96b90215cd7a170d88a42b53275cb49e",
      x"cb4602e8c09dd59fc2e6dc65bae8c849",
      x"8aa6eb5c0641dbd2fffe61dbaf4cbede",
      x"8ad269a1d26132864bc085b0bbeb1dc7",
      x"fa872700bf4e227e127b8b5eab61445b",
      x"026a0fcd87d925cbe6b229e38753e3e9",
      x"6548e2cd4aada59c6a00ebac06d342d9",
      x"ec96dda9184a22ef9f965f16f6eea039",
      x"397f58124beb92021c91ba96f897c564",
      x"b3336d000aacea0a8d3feb02c443e27e",
      x"03d55db43d653378176f2a9517e3bdc7",
      x"d97636960b197e12ff45eee71eab8cf1",
      x"7f6afa34daa96ee91108b1d613fe0dc8",
      x"bb9b240fe97001c51bcec49263c16b78",
      x"ce736efaea748a0183c04e4698108464",
      x"b22d36df164236731799c2f154d2fe9c",
      x"cb6d5c81ccfecbc62a2277266873b030",
      x"f2c7e8fcb8288c835eb1857fe2150b4f",
      x"772a7f35934d569ef4b44f271e420bc8"
    ),
    (
      x"683f6478b263b6df257f67a44eebe296",
      x"168e2195c8ac90c203c95ebbd7b92803",
      x"5ddf08bfeb8511cd5807057c5b19078c",
      x"648fabed53712496e63295e39b060d23",
      x"2186d2ff74daea46d7c2b84d47bd732d",
      x"467727e023e7babf087f2cd7364dd4cd",
      x"7f4ec44132a6da97dcc28d9d71794c5f",
      x"b3818daae8a76a522b8cee68b3df5c16",
      x"585b5d2fd7e4d3079834a2ab9d0f2a48",
      x"a3a06ec87da0774095ddefc06d72182d",
      x"de6eee1dc27156d0be95becc913e346d",
      x"00028ddb25d316c29017983fb4925410",
      x"5c2f4b9ff9749b7e445395e36768f6b0",
      x"bf3936e7f70b903fea635745109f6e5e",
      x"c2ef460f65d8edb1a46cb24ed89f65ee",
      x"d4d0b779ff441a9e272293e3f241baf4",
      x"c8b70969ae36a41ac8d4bb23194d893d",
      x"e8ad0d6fcc365d83db9338a60ca1f592",
      x"23f20ab7f70ae73c94d39c57dc3b332a",
      x"863e4c41be196d47be9818dfe0f62f91",
      x"fe71b032e634146bde3d8f63f2dbedf9",
      x"893b07159416c400f60f8e6faabbd2a6",
      x"646d363743e559b96b2f7043ea197aa3",
      x"f1c92bcd47cef88957cd370ecca15ddf",
      x"18d5866571c46bf32f7e8d4bbfd95365",
      x"34d13f9441af09b7dfcdaef45f7a8efe",
      x"a6aabf25e8854d060a9acc3a69d0fe70",
      x"50262be21f9fcf0c0453e988f30fa00e",
      x"125c9d7cf069060fbae019204e5a1e14",
      x"a43702fbe370963ef36c75d8a8b6cf2a"
    ),
    (
      x"676633d87c8c6781c10bc25ae6f75878",
      x"5961adb11b7d30ee7b499fbb41b7b4e2",
      x"47c338e1beb9d93482d31165cac78547",
      x"cae832b4d2388495a528fa2901cf47f5",
      x"40913daf1d44bc32d04fc0e6241a0d18",
      x"8e1aaad8dcfab9029249a362e0c3afc0",
      x"7e1b96b1bce08be5d4efc5944ed90ba3",
      x"fd13db9add8496b80c8e638f8d4f06e0",
      x"7ea9f66a4364d87c82aab648d0c8e2ba",
      x"4a9afaad839c4a8090cdaa9febdbb639",
      x"7a8c0d2dc3dd4a9d6dd7d1074004344f",
      x"3fb9bdb9ef52c1ba91153e3e5800bbd5",
      x"b966f449ecfafdedb5e2c2b71c379d4c",
      x"da4d6c1ff47740838b4ba600d8ecbed4",
      x"4e78424f70bb720243feb33e7d4c59ac",
      x"eeb24eb6343a0410b832eb620b3dd2fa",
      x"011532ee86336424642ee378e4fdf774",
      x"2adb2af983da0ff53c2e3f7b8a5b22ce",
      x"4ea8bb5c8bf2d397f44cf95ea0f480d7",
      x"4adf8dd9eb1ad7032b05f9915fe8dc11",
      x"606fe2b6ed3a07eb5f362583e9e71ed9",
      x"eadaed902f07b1dc74439183dd3171f6",
      x"35960075bbe87f3d521651da1146880a",
      x"09a6db7547749ec9de5b221e6ceefa72",
      x"d086c33a539a369fbf087e4da5ec73a8",
      x"71746feaeeebb86f797647ebb947a40a",
      x"6e0ce5d8493c49ff213407b32b81692c",
      x"98974bf6aeb99a0cef6e0db4da4adcf6",
      x"8bc507139b7e2b8b1cb484e61c7cfaa1",
      x"9af75b7e1a9fb3de1a4d4352ccf30449"
    ),
    (
      x"85ffe3eec111c19d8a8f7577d17ce43d",
      x"66e6cfba729a12846fb186ba7da1942a",
      x"6b01282ae106097a7e090f7cf0672698",
      x"06984683c10975970d70ead0e1bc6f8f",
      x"bfced29f488f8b6b448a1e7006c2691e",
      x"8afce995bd7863829c1152c982f35e3d",
      x"6e2de74db0a626c5aaf91a76c512086f",
      x"c3f953049cac9c0fe32805dd9776dabe",
      x"bbab7b68998e4f02b2fe33f56f2a81e7",
      x"1841daacd7acfd1720d1b5fd36f0c18d",
      x"1a63c8a88c3e326e2e1de0520f9159fa",
      x"cc84e6d994e8b634a7f9d8b4ec0e9a01",
      x"d262ad074530b1284c68e99a913454f8",
      x"5c289b25059af1a79839e90cef4eb7a4",
      x"dbb4c22b380a05e8d800953fe41909ea",
      x"cea3f3bb9e79b03b491374d6b207a15c",
      x"f3f2f20ac8328ea1bdaae36ccb060d02",
      x"492fba54ed1675769b063c17802d36cc",
      x"94557cb30b4886d38ccccaebbebc7b78",
      x"a98bb62cadf4abc40b8123ede9382459",
      x"7769005101ee7df0fb6decf425d74cde",
      x"7f6cd22bb861526abe6dbad97d42cf73",
      x"878c0e05e0a6861d52a095fe1b1260fc",
      x"cc05a0290f48e38afc285b0bd49b6082",
      x"b086ce239af16b1c993a71a872a4417d",
      x"ddeb7edb5059177136d3c26be63d39c3",
      x"3c7ca7b05abb1444672a8dfd7fab05cb",
      x"dedafc271a9e2574590d388edfb5ab94",
      x"d6b924a0fbcc4fa8a3a3014b25adc5c9",
      x"83d1d027d4c4908ec53ac8eb132cc8bb"
    ),
    (
      x"449ce29accc0eb8bf13d17deafefa5a4",
      x"99e888e308903ee8bd13f0f4d8f026b2",
      x"0e29cb2fe7ec6fa9529a23ebc6cd8831",
      x"3c5957c28db246e62e1758f93e9d549e",
      x"e845863834f668a55bbaaa101d21db3f",
      x"c8278b3b3aa22640c6291ef5fe387080",
      x"34e896e0dbf1a6a34acc2781968354a5",
      x"a7e27de05a0a532ddde2b5736705ac4c",
      x"ccb56ff2d2ca3219b2614b1e82597110",
      x"14a50070b9213830ff3377fb893b4bee",
      x"ce1f0b58a60eccf549f283d223cb319a",
      x"b10efd992fc51878c3b8e2adb6e73ad5",
      x"3e99b351469731df2a105026a6fac996",
      x"5227bcc5f433ba93e2c5aeef63f3a592",
      x"4396817c6f0fa9a3668d0ecbf5fdb775",
      x"9d0a4d4fabeafaa10f923065ff654c70",
      x"53a48b9c65200320d49e18366ef66cbf",
      x"3d35d5db79f98287285aa0af62e84ae9",
      x"55c585b2c7a2a5b6a4e6f3930a059843",
      x"4fbf4ac2865e533d9146f8e9d51d216a",
      x"55486de363c79cbd74c42201115d4bf2",
      x"94940ec1b821ee1857f9293548ed015c",
      x"a08cb63c02fd54387cba04ba63b1c372",
      x"28c6bad1b70802b5423abd8352bad8c0",
      x"2aafb420d62b3c702685734ad12bcd60",
      x"1b002a38f85fadc93be1d8d9226f99fe",
      x"847b57ceac965db4e559cb0e796c03e2",
      x"eb0b2a499f0f98383317b4c7dc616cef",
      x"4668fd1d6844fa9037cbbf5dcdaa1e7d",
      x"54a73d0ffc109e1c03841a7b55738223"
    ),
    (
      x"0d47faf7b2af1211ae4584a1b2d2a91f",
      x"98788e38a72eca1c4e37237235e99c89",
      x"a8c9e5809a397ace898de4d285ac0637",
      x"75defb7a31e1896fa78573cf783b76e0",
      x"6a1e740a8472403f356c94fb0f41c794",
      x"5bd573aa1949817778e01076bc8a2028",
      x"8e979149fe363209caf37e2fa3fd9624",
      x"aba32fe9e798551cddb3c7170191c649",
      x"2d93d956e2250c2006431c6af843ef72",
      x"5c3fcd7ef6fa8851ded39339e966a6d0",
      x"ab91b30ba805716936fa62e4879aaae2",
      x"bbbf436d2e7c1e4080399f939e61f5bd",
      x"8d32fd7641f3db00beeb29cccacef18c",
      x"37ef9b42970437369daceca751f10be3",
      x"164ad08a02ac78096e96b74a2f55dd29",
      x"244129305e7974a1401fd8b6a87bfd8a",
      x"97c09f5128dc6b04f410f5b467f3a3f1",
      x"2c6d256dab04ece3ea96fb79d598ff81",
      x"00480be984b753451e2683ab4780500d",
      x"58868a38670ff47fd01cc8440a0d246e",
      x"a57ec1bccc2ca906e15ccbba8866a51d",
      x"917ed8c9f7ea81cb410b75ac3d99bdd3",
      x"ed3f6cf73d257ca2fae9421bdff76d9f",
      x"774fb680a06f212ca0c27f1c32111002",
      x"4332c28d533cc394e07cb3226b4b7a7f",
      x"e0ef58acce720db2551bc82791dc9487",
      x"6e8da7c7ae993aede359c9c7d7fa7236",
      x"1a9384fc027d2d38a08b3a44e3d957c9",
      x"b65f58573705711266789d9aec296846",
      x"cebf85a3a9b275fc807aebc0ad5cd845"
    ),
    (
      x"128e9f75e67563bf05cffd1503d8680b",
      x"01deea243bfde1933342b3b905c50e0d",
      x"ae22187fdd9fbcc2826e3da4fea18648",
      x"23b19d43364ba21b855934b0ad9cd677",
      x"00dc46e0f78706c514772e48593ee170",
      x"7ebad13f93555203818d9e0c0c9e2f29",
      x"6149454b4d317f3d368b2e8f18113686",
      x"dbacc37e44d9116af9bc0aa95f72e0f9",
      x"e9df559c426faaf943068368b61cc1ff",
      x"a49fcb21a3285473d94f4574d3762f71",
      x"90df0ae68ade01368048ed6b6099f380",
      x"f94f93e7bc214c580086efca1032a373",
      x"7438863db3eb4a8a059d1a02da6d7a52",
      x"d1ea25e580b8e721c2d64c58a1188067",
      x"f14663e6bbaefdd609a790e0c20a06f7",
      x"41a10d8a0134e51ffb7d214eadb194a8",
      x"ac177475bf86051dd2643dcb87c49ffc",
      x"9527c3d03877b3e52f9eb3d18f256f9b",
      x"6b454f03e068478fe3e3147813353160",
      x"c280dcca219ffeee538f47a2f307ba63",
      x"01b99f897421a8ebacf7319a438a9d75",
      x"748a93c7ee6605098ebea3aa00d7ff8a",
      x"7edfe9a9b43370d02a626885a4abe407",
      x"2a003dd8141ff6e2b4a94b259ae92141",
      x"1a8169dda632aff2db76c429d0e4047e",
      x"559ea5b6e8145aa865f8fcbdc2d17dad",
      x"5276951bcae5a2bc77bdab11926de924",
      x"cd20993cbb7e8393593a08d2e3b18a7b",
      x"8a74f20c78f64ef44809f6a2a19e110e",
      x"42270a584a9d92f6ca0798e5300537b9"
    ),
    (
      x"030e0e8c5d01d887df1e3885e368a2c4",
      x"51adc6cb7b5d561650dbf58ceddcae16",
      x"0d7eced06682ac652f77b8c235257e13",
      x"4dfa3e6701bedb30a24209605b15e67e",
      x"9ad525dfb762d4074938a703432064ed",
      x"de1e4050f2e81a44f2a5d2cbb95536b9",
      x"ee79dc25d261c5aec1810ef9055ece57",
      x"9b74e2daef8428e968a72f781766dab3",
      x"a4ef2ef91b1b7940452ec3cf2470bbfd",
      x"a13870210526041a3a6478ad9365e35c",
      x"b08b878a2b6497a0c93bba3d0d44ea22",
      x"d567077fca7e7ab4ac367e900b8cb4d0",
      x"b223471f1f7f2c84a4753bcc34cf595f",
      x"8464e8369db8b290740bc5fa2ced05bb",
      x"e4cf3f741310d71c1e3bfdd36fb4e9e5",
      x"ccd1520fcf3b1619612b20d1bd57fa2b",
      x"51b19285ab8da25bc438a4a96ee97fbe",
      x"c06b0d57d8b7fd0aa5d598f68e146233",
      x"5e7670a7759c5940b9870f3566317fcd",
      x"a22db34d974c3297ac197b42529709a7",
      x"a4da2525327a0618a4a1b5b6b863dec8",
      x"021b5e631c6de7f89dae3792de842f2e",
      x"b7b3b6bc827e8d6e891e5f47d63464b4",
      x"3adc5eeaba21a35901a8b57f0c96cc5b",
      x"36f37c97490bcb3d27cf12c44f23ae6b",
      x"752d00bafccdd9490e8082aa5c818607",
      x"9758ab867851e2808e2d3fda80c17cba",
      x"d72a517ce79f2a0eca7e3c03ccb3d10c",
      x"f3f7334c0f525d9d8ea1d2e1d47f6b54",
      x"a912fd79c578bfaf886813e527c861bd"
    ),
    (
      x"26487ce0601d87e879df70f872745983",
      x"2b7cc61a172b909f2fb60e2eb312c42a",
      x"078c438e1b7ced0c058554f77d7ac9f0",
      x"2eb2063adfb98cb6a78e965eb7a9436e",
      x"ba30f90f4457f84a73767de55a188779",
      x"0e029c7b8b62d8fea3febe0ef3ac1877",
      x"a67a5e120213743303e584e55d6991ea",
      x"e944f09ab34d4ff6338272d7f487b368",
      x"e0155e0480fc78982f6a301e6b8da3b2",
      x"5d0d648ef30a381c5dae8c7e0bf13935",
      x"8f235d72af062ef57cb2d9477fe8825e",
      x"438604cefeaabcbc6529de486b44d0a2",
      x"eadf3bbb85ece44c94e57b412b982e15",
      x"26d61367014d044f6fd1e7ed9126a19e",
      x"ab8098a2fa23fe5116352ce7354f48f0",
      x"902281b67390b7c4c2042cbc2c2ee165",
      x"95c309f0bb16c18a01c3d0e50f525080",
      x"d276042ffe7af1726bce1325975fbc3f",
      x"168819c1cb7d2bf3260964bcf5892e03",
      x"c88478fd88cf9ce8b69462a8a4052b38",
      x"7950b7ec1a52270d9ffca00728343e47",
      x"43aedd5391d0a5674812a7d400f62871",
      x"348cd20f256515f33c9b06aac253605d",
      x"ca12c00512c91f4717d734ed852dd7fe",
      x"5279a1adaf93f8be1dcd3bbdf60782bd",
      x"6b329dc647f664bdf9eee11e9516795b",
      x"e8a12f9a7577b77c1cbcb4c40b1cc9bf",
      x"2941b4a9e8379ccb68ebb032bb7266ed",
      x"9b68f868751338ec0358e99764febabd",
      x"da9a807ef33e6b76abf079027f508695"
    ),
    (
      x"4a7f57ba225d641cc91f708b72df7e0b",
      x"b17a2f9591db9caf6d6d75f8825c935c",
      x"01931fd97ca3791b3dd2bbbacb62b150",
      x"fb442e9b482fbaecec26e42d622ef8ac",
      x"048ee142191e2d2b75cc5df4f49668c1",
      x"20583a036d1887d0c3e798fccea05f02",
      x"ea4284f911ba01178a8bc5964a608b87",
      x"150749abb616e28f3161c9cbb0c8b3ae",
      x"2c0978b1e8f77dc5e02eb740c0f51bf3",
      x"81ad9ad1c51f0bdf0f062db55b8f5926",
      x"70b7b707423d777558c59b514054462e",
      x"db124378730b04946ce94d3533fb9fbd",
      x"47f9bd6476e0901128304294dc6a6825",
      x"e00b57603a6276a5c6277789089675ea",
      x"4c318f138d79e40ced3990389ddf485c",
      x"571c1487d87166f6faa3544cdd8b086d",
      x"70c989815a3d23d0a6dd9eb60c2d48f3",
      x"f5a59d02611e350c28436a04ee00389b",
      x"a9a0e4c88abc80c12e4a1f7140536cbc",
      x"6ea79ba7ac2e17d02374285c0a3a8582",
      x"e23033749464d60449b9f98bb0ee4565",
      x"a9d79b51ff39993a3ca4f5ff99bbe0e4",
      x"d8a3ba459c7a8aad2bfaeb275da29757",
      x"532b3f3093ea93fdabddb0212e2f18e0",
      x"80f5e40870d9c4a2c4debeba2109f8cd",
      x"be8488bfb46b5d7b51257eff7c2b0de6",
      x"7eb8161640ebea73dd276fd51113fa3a",
      x"2ec5fc7e497e830df0f11aa83c671377",
      x"20deac4a6f20de29a29b438b0940f440",
      x"1c31e52e908ca3af9873592e7e713123"
    ),
    (
      x"5e7541e9aea84b411038e8c941d415c2",
      x"4b355124d22536866b2539766db68c12",
      x"4ef71a79f4e1e60f90aed39d51af5d43",
      x"7ee98ea072687dfa1485205906ef7ea8",
      x"743afe57779b276be8058a867d49aaaf",
      x"a4660096425d5b7ebeb648741e471bb8",
      x"95f32e30848bb9fb5ee93a83f597db33",
      x"58d4d61482dc80aa7203d2eecdc7aac7",
      x"2167923c8d8541caa032ec0493de97af",
      x"5723d5178c072f87bae72fc898f4b0dc",
      x"d94d3620786ec17254ca650e816066f2",
      x"33ce113aeb35606a4bb6064a9b352b45",
      x"f3a0d1f41cc6393a807e59e99bf15758",
      x"b3bffbfb9b90529dd339f91937d93517",
      x"6242f6ad0c18173be80324f6ed0f8f92",
      x"26ceacc1bd5643b70a81e1a4bb141a18",
      x"80eb232e43de5f4722f3a2f05a74575d",
      x"e29420e773707483414eeacc0ae9b6dd",
      x"2ecf96b1aac8288776105ec5699c200f",
      x"767526c1c029ada057c6a3a0855edac5",
      x"bc4be4f6cdd1f77bf6494f8bf5246542",
      x"db22e0ae80fe29cf5ec50a6591242f63",
      x"cf1df75e32f760b3138686855ea83103",
      x"0aaa673fbbfca4ccecebc8c9c77e67fb",
      x"9aec755db7aed424d4c5876789b7dabd",
      x"5c86a00fbc4883691fc5fd8ab6714f76",
      x"45e028b77286095f347659f0c33f5f9a",
      x"ee803801dc40fdb33bef6bb45aa93146",
      x"42e0268c41ca18f5ea07ff3015051285",
      x"6e7ab42108015712c23a314b63c4c2f8"
    ),
    (
      x"b59c2fbfe36be28fcab0e989cfe84315",
      x"d060647636a0ff9400a70ca3436a852a",
      x"b445fda3d4a2ae790da9a30d6844ec15",
      x"03a73ea5b2c4539205c326d3583d3e9b",
      x"4ae7259cdc6af65db1d1ff1765805098",
      x"71970f21ff28622564ad79820ae62ad1",
      x"8c6937bc82dfeac6f6e4ee55fb73e5a4",
      x"3fd9cf593116549e045514e41c004aa8",
      x"605c9342e69fed2baf390f3006671bf9",
      x"5d74697451b414d7f27f33adb8078300",
      x"172aba03abff8b07c4e9982ff696a821",
      x"cedb12025f4bfe03ec597240d469ff98",
      x"26a1aa6c4a02c1baf35bdaefb50d7dce",
      x"00bfd974e8e1497f6934cb46c80fc693",
      x"09b568c770b49781be1383570330ec26",
      x"0de7bc3dac27fffa171ecefca24effa0",
      x"39eb1a2e122fdf3a3f167d112d7b8fcc",
      x"9c85b9c3861d2850bdd2c88ee4286b53",
      x"14df7309389ec311f3825f0c8b5e5b08",
      x"f39e8232dcd94ff5c284106667fc3106",
      x"721cf62bc47e2b3cd5f075848df89248",
      x"6e48327fdf7c372b7b737f832210e3d9",
      x"97557d07cd0e74800cd1d379f0f8d05f",
      x"7d261f421371a375d5f28930510cd4d8",
      x"35aeb085d9470de9d72d7d640ac99a5a",
      x"bffb8f674a96bbe8c61b5c09249dcee6",
      x"115fa96ea4ca4809ce6fa86e78268241",
      x"d5b84e7fe738edc81d1eb1614b945b7e",
      x"1d6698603b50562c35cbf12dff2b91ef",
      x"80b2968910889aa0489e7dbee7d01d8e"
    ),
    (
      x"bec1540d39a9c80c1e7fcd1a7310b39d",
      x"9fa383df3e4bc61b1bc24f6e32cea283",
      x"563350313e7e6753c7aa79b916bbf8f0",
      x"2c7e6136b2fc1aef53407f15295dfbf1",
      x"be9a67a809421884a9ddad24fe494f64",
      x"f8bf39c32522ce508c9175ce2cf2e269",
      x"b0b12514c04d082703fa1b7e2932bf78",
      x"600c49968dc3894585508076613ecaab",
      x"3a703a496a4190dd5c50ab645afaa80a",
      x"174155a5cabc7d8a270e0e87639b7d9b",
      x"a5fd1cef69af0f2a17edc47f5900dad6",
      x"3ef01ccdd474281e4a9332d4b4bdab80",
      x"78f836a628dba5cd272cec4432fe9309",
      x"50eb2f21f18671676fba623fd51f4f1b",
      x"2e31b3528be10f809afd3c58fe0ca4fa",
      x"e059dd23d48b60b28a4e7a9ec30806c0",
      x"44ca9da75aa76d85b3872327770ac54c",
      x"ffcae2c51c8b01e95315b1ea51bfbfdd",
      x"c4443b2a53d1befc25d6e8dec60a5c3d",
      x"2c69f869fa8c63b35a0b0b8a567426b4",
      x"5feaf433819b8e998ce3dc8416558054",
      x"6d3af8aa558e2e3155139769bf76bf9a",
      x"33a1eb81b41aa5fd699a6fdded655116",
      x"1e3ede616859792803e9f018882e9aeb",
      x"7570123a389c46c7db3e67d6bc684d39",
      x"f3e0585461af168aace299ed84cb0a1d",
      x"766d3f86f01ff0b9372b30a8ce1d17ca",
      x"232455e5af116aaa83d6aada3c751ff6",
      x"5ad0f942af87ca9c5184c73a7ba58729",
      x"ab6878aa946f5d3ca772ce6ea2d00994"
    ),
    (
      x"83f432ef1d3593287c73d18973c733b5",
      x"1b7e10067cf68ac0ff4c1abb3c202ef5",
      x"d431d32356141ad0a24d9e1958a2c816",
      x"de43624b6bf9326a47ffc656d0409ecb",
      x"d922024d66d53190198d5290efd6bf75",
      x"066d7b099186d74643cf8de5eebcfda7",
      x"3950da988336bcaa50fb10137a1a9407",
      x"1e7a4576f7a8bc2d25f6547383aeab33",
      x"cc7a46f49b0ec8b1a8c3b32257f742c2",
      x"0e0632c89796177ba33d1c14223b824e",
      x"98a35d0f1688f006435e225998b01a2f",
      x"e04ac3bef76d672590f1ee494193c4f4",
      x"6f78b8acf703dfc3ca93c04cfab7f119",
      x"9831ab3952fc42bb5bf8b08fc9d7d14a",
      x"f5de75a58920832f8709d03627a8a722",
      x"52455f3d22f4f2a471ef9c8e4ce10d4a",
      x"69055ad9a0c57ee22f3e39307b5a48a2",
      x"7bc913819c6c20871679b33471df7005",
      x"320a5b2a23e2848e00502cd6737a559e",
      x"d5660043f3ecaf1bfa6003b5f2f75033",
      x"27891bbaa1d970b9a36c969fc35e1de3",
      x"5790aa75a0034cf418d686e7054502fa",
      x"baaad026113d575921114b8c54b77f28",
      x"219b403f4b4cc26838506a2bd6b5e91b",
      x"81bacaa30b7df93cd9fb9b70c3131019",
      x"38ae1a11fb2d615807bbceabe9d59c1c",
      x"bcc6f3dc9ed54c3b12c3ce3f9c6999d8",
      x"c8ea41e46e7a0c6822daa976feec21a1",
      x"a7e694a0f04b84059ad4ce657af02a7d",
      x"e0db4dc12df6f864d083983c03e41fe0"
    ),
    (
      x"954bafb8292601de797f53517e3a450e",
      x"823ed3dbf29c64d420ce4b9e3df0fe15",
      x"38bf5a299ece2bde222a884d0206e0e4",
      x"ca8215d65dfc082ed9924c863b459a17",
      x"c2e1cab648539fe19452173c0394f9cb",
      x"c6e38a87178b357e4242d308c500f582",
      x"b0fe92382facd84b30245e762c52b6b2",
      x"0dcef2a0dfd4c014c98ae60b7a9d7d5b",
      x"e294158327ca21d6fc10679040dde44b",
      x"b2ac5db5183a9a9fc7b5499db9f97a27",
      x"b2764d70047157f5eef4e6548141e2c2",
      x"bb487eebd2ccce79983474bc74064bae",
      x"460d02a2be3863b35d12eb8fbd513567",
      x"54c3427deba5bfc0f067395b67760f95",
      x"fae961af0eab18c77a60d53d931bc5c8",
      x"9e3461fa86bdbcbecbfa72273c9ced09",
      x"ee266754998db7fb8804b2ae9fa13d18",
      x"be7eaad6b25cf97f758004e76fddc68b",
      x"3123660579582397c2a16f928433a636",
      x"f7950802a1dc4539c9c66a44d03c69e1",
      x"c1aea156d1f21b2aea5e25a391526073",
      x"90939d728f4c9d0e92a35f1cb28f51de",
      x"bf63cf616ebab4006080b82e38a01c56",
      x"e5169db7b0cab99c81a5ecdbf796220c",
      x"ba8bbc1c49d64585d721728acd2231b3",
      x"e4ddaf1b7aa5fad1762cba11a6d32f9c",
      x"bfea3d61f580a16a4b5dd2c75d8f4b4b",
      x"e11013d2794c7f750fe3b7ea2b5286a7",
      x"59adea0a3a653dbf8691b253c602ecaf",
      x"06316d436a54cf82d3eec1f15d544421"
    ),
    (
      x"6deb1a3c6045ffb01c2e1dd8ec8d0fe2",
      x"1f0fe236625fb12712463822b2629610",
      x"87e63a7ed481460e5b98b405442d9707",
      x"4abe6f2d34cde592f23a2819b583a033",
      x"5cd1d3e5e5d1902de5b00d9ff9541b48",
      x"0d8de3edba335707ff65154d7008ed3c",
      x"c1542b357e3b3d5602c38078862025c9",
      x"585380acfa0e378b4e6884671feb0d1e",
      x"6f2f0c720a4ad62a36d7d31f601e29e4",
      x"263da3f58f0a85147d588b49191fb837",
      x"be82eb31f608befdffe3411962d30d34",
      x"254f6f9c9f7d830fb0701cd6c70001b7",
      x"46704d7c1c1f1a759491758bb27341c1",
      x"3ef4b134c57e23fd1d7fb0e61a4da01f",
      x"4e371a6f96de0b29e270c529f8fb969f",
      x"e2b85b03ca15171e0392514693c6382a",
      x"1a085cc6255a1b6a2dcd9e3b0b87dba4",
      x"36facceb38a5a906711e333198da5091",
      x"613147e1add31b2dcae45881da3e134a",
      x"43d3ae11a79d69a42b808b705ee46e67",
      x"724ec048942cbdadef6358c0f81e7015",
      x"1bf63e6503bb30c3dd4b5de0950be08a",
      x"2eb1549080ce1647c1546b5575a334aa",
      x"d892fe95d1c68401c888bb423de10317",
      x"0176a6d8166386cf50c97151ae69a406",
      x"75776f9e4192fa204702256ac4a73b71",
      x"74b20fd3cb52af64b5bdeb5a2c8ac130",
      x"2e625c1f88ea8634a4f1b4fda6def461",
      x"7306dabf2df3cd5e417a5f72f02e9331",
      x"90de0ae2c967a2ef0068a8c7425394cf"
    ),
    (
      x"d8ccfeb0068102f477d0622467208b7e",
      x"5b4538be311e2bb37f3e7cedbe4bb61f",
      x"323634aba39ee77e17a2efced7f3f31c",
      x"556c605daf51b792f8761e8962f6345f",
      x"4ef0e9993f60cc75544f7a16abf70e57",
      x"8cacefd2d34c34a88390fd049a02319b",
      x"f40ca5b93250da86633d8d528dbb8a78",
      x"a07066528676fa246c3f6d2a73f11a27",
      x"d6f7a19cefe60001181fe75de2f02ed5",
      x"b412de6f0872696b33e8110ce8bbe423",
      x"3b4cc927b50a66da66660d7ea0195031",
      x"3817e62cda9a0fab59b37f8688b6b011",
      x"7bcabed77728e78e662c8002b3fbb867",
      x"dd4d78538f15d17c3e63aba56c2b9601",
      x"646d0ea70e2aec8421130d6fcbb31e68",
      x"5a9f19ff933f0d8a722d76036affec7d",
      x"37fcd297d411cf84dd356cc1849c235b",
      x"5c64999cea55f1f8d6dd98cf0e7176bd",
      x"10792f34cd1f968dceb0da2f8202a141",
      x"824a5cccf865ea7ac9c9160171696c3b",
      x"dac3b3afa204c32568d5853f112c1c55",
      x"ccbe818cf0f555475c56436e38c0b0c4",
      x"27a77047bcb7b5e9958195977433a56a",
      x"d6e24dd4cc39705bd7a7c6e16a5ed97a",
      x"a2f0d58d479eb3c032dbc9738e69cc12",
      x"4b352516af0a2fef9025b458537df846",
      x"247c79a48f9c447726b1dae46aa4ec80",
      x"26e89d053357364f665b9dcf037519f1",
      x"fe5ff822b9a9f6ee72119a2c930bfbd6",
      x"73423df0824991a3571aa6ae42385eab"
    ),
    (
      x"6e71275c3920c5237a6d4a2ab5dbe92e",
      x"732e78a0f4296e9bb3eea2f44ab6fdf0",
      x"066df291982e1fc0e5554c4ced0686da",
      x"2365e1f227e7b4af0e566726cce047b7",
      x"ea888667aca04d9064db997c23c8df3d",
      x"e90c3b58671e8d58ef38fafaebebdac8",
      x"a41aba2831dd14029c23591489ed8c4a",
      x"23abfbbb1ee87f7fae3694d85acd5b29",
      x"91f5dc37795934c59a36861d7a0e08c5",
      x"679c6011cb5e66bd4b6d0a25ac8a65c5",
      x"1acd97fa5b05343ae3bd6df95919e857",
      x"2cb1b66f4f87af656be708081bd37804",
      x"0a0ef95a6c040a09813042fb69d1356e",
      x"8c1d14a35aa823aeba93416419039c12",
      x"065193d1130273d07aa29f5c398748a5",
      x"d88e71a20055ee861eecb5f5e316f270",
      x"93438ab61749010b8d35a1b0962fad50",
      x"a5ed560524b23db74f2291610b5c111c",
      x"7db89a5aeeda13c90cf5760be506023e",
      x"205bfa1760ffce282e7fd1ee528052be",
      x"f5928dae61df732a26a69014597930d8",
      x"ea1890a701b31dfaab23763d0bd987a0",
      x"871c6ebc151184e9c7a59ffa3f461de0",
      x"cf69f6dca1d1aed0e3f4002c1851ea9f",
      x"b2214dd8740cc4dacb8107596cf9041d",
      x"e22f92bd4e84a6e2bed3c084c4e6444e",
      x"83c498c905c3c6732ba8a5e8af8d9c33",
      x"b447f9383cbc2491919cd5f3a05d2dba",
      x"511d44535a1469e20d010cb226ac908f",
      x"6e875316331ef5bc80ddc0817632c7fb"
    ),
    (
      x"f5ab0ebb7bb8118d349f5732ec57f5d6",
      x"bfb4d2482e2ac38f22e7f0ce894b0d93",
      x"fb460334d675d210e2fe16b55f284522",
      x"e08077cd2403138af9dfb1647b90e3ed",
      x"2bb4e2061a477e54dd630b014cce23cf",
      x"10e36f12cce8f189d894c1f36f6c11fc",
      x"6204c6a8454b35812d18ee04cddff292",
      x"2cd6b38b97e5a65751943339d6b0c4da",
      x"8f89cef5d6b06d3fe440fdedc217e23e",
      x"0786b34d75a9ea6b89934337f69bb119",
      x"b15600b44bf364369cb1cb54764452b8",
      x"f89ca2bca384ef3fc530bdbb3e01b4ff",
      x"5a83878197ead0f42f6b7f52ed38d460",
      x"d035a4ef987c2e60e0a85c6ea6f6f217",
      x"26b738dbf608833df52a529791d8bd09",
      x"a2d79741ad667174f1ea91ef9c5329b2",
      x"0c8b2c96a3bc61cd7b88d8bc4d13feb4",
      x"0a68eabda6b52707723641bcaba36425",
      x"4fb0e95bc605633533d6c421561a1468",
      x"25f20dd61b6d6c692d0afd5b7e5108ef",
      x"91b925f053654a09a6e2edbc2a7a358a",
      x"1df628162dc27f7d1637549ccd148c36",
      x"754daf1c4969236beb44d595f6f88d59",
      x"d1927054facdc89008f9f0c27f2aafc9",
      x"742e6e2d8d0f66003ce250f8671eed74",
      x"c36271c2d3cff234408b7fd6e457ad87",
      x"35da472f2081a41a8c8c6240de5bc2df",
      x"821dcf20d0f375b2e562999e7a341466",
      x"d821f67f9cb271e1de1555afa8254afa",
      x"95cb93cd5a0ee3413942383f4edbd855"
    ),
    (
      x"d16c343c9f141a870021de9149a03475",
      x"3f6b0e938582dc9f3bf528b0c7213e6a",
      x"526cb22992ec1cc67124a329d12ada76",
      x"e7d65a29ef9974409c6dba3ed5837745",
      x"a90ce717ab7e6c419037232a5817663c",
      x"ad9775af28daa9059be4d66161be05fe",
      x"d45bc3cfa9ed6e8e0066341873266a90",
      x"84afabf6462cdecbaa34aa9dbdd7e1d8",
      x"c64d695980aceca22a2f81a459a45bf7",
      x"d21579da38bd51e7819a68df6fd72df0",
      x"8e8ad6e9cb72e8c7042baa038843d1f2",
      x"040897015b6abd01fb68456ea191a7ae",
      x"f2b41fb5c1906623bc08e26cd0e913ee",
      x"da3ce3aba51c9142cbd0ff30263b6c8c",
      x"0f272cd2104043c9bd9a6b7bab839b45",
      x"4506061266cef9adadd9dfb89d92331c",
      x"60e78e5042b7f9fcb552280ce3c61e5f",
      x"251f53e57d416a0cf86633ffbd890e82",
      x"aaf34b97fb9a98ec948956d0b7990c54",
      x"d13b8fa06f1d1f4a97fec912d1d80602",
      x"49366518e411fdeaa9808041ec083261",
      x"d7ecb020d9cd9d5d8e3db66941877d6d",
      x"e4a941dfc10d8886e50506d503332939",
      x"75a343449555c3f58ecf43fe2869046b",
      x"d3a95bd293628d8de01e595e417e5f58",
      x"48790bfb7c534fc02ce865de89c9cb58",
      x"59ed2e74b64a5419de209acd0fc0b386",
      x"f22dda92be29faed5b9528d2c38fc851",
      x"9c169c9450579868ae5d077e1bb156d1",
      x"16e8de5576ec038ea97166b4385c9147"
    )
  );

  constant C0 : std_logic_vector(N - 1 downto 0) := (
      x"000000016ee016559278ab60a47f1a8e"
  );

  constant CONSTANTS : T_RS_MATRIX := (
      "000011000001111010101010111011",
      "111100100000001000101100000111",
      "100000001111011001110111001011",
      "010010001011001000001100001111",
      "000101000011101101111110010101",
      "111110001100110111000001100101",
      "010011010111100111101001111010",
      "010011100111101010001110100000",
      "111101101001110110111110101101",
      "011000001110110011010100010000",
      "011111100110110001000010000110",
      "001011100111100101011001010011",
      "100110100010000100101010000001",
      "111110010001100111101110000001",
      "000000011011101011000000001101",
      "110111101100101110011011011100",
      "010111110000110011000010111010",
      "110010000011001101001010010100",
      "101011111100101110001101110011",
      "010001111101100101001001011000"
  );

  constant ZMATRIX : T_ZMATRIX := (
    (
      x"1937dfa54e4c9940921f3c5421796692",
      x"34db8057ab9cf82bd4201f4d77dfc788",
      x"28ccbc181802fcd6a04bee0bf11d1092",
      x"8370019947a81d267cf8dcd8dbe40498",
      x"c55678c0770419d7085a4db47c2e8282",
      x"ef273e4ff9afccf13c5d33c7b870e7c1",
      x"e56f68f22b4b3d7755072f3c7634e841",
      x"c3d0839a423beba0c868ae2445a00064",
      x"1502ef5810a21d3f29f50cb19a871365",
      x"cbaddb72abc93466e8195df8e2be5d46",
      x"5d2929dddeeecf48e81306aadec65d52",
      x"5ca1943cd287a8174d38acfc4be8c316",
      x"847901ef1b054de6553eed6a7c794f69",
      x"842b2f82e9bffaae19a5f1fe50b04f17",
      x"5011e94850b95937adb713e74e484eb0",
      x"d43b055f152beb2280ea1bca1590268f",
      x"40060c1b4a981341d743dd1769840799",
      x"975e5a3b184ae8b6c243df5f873209c5",
      x"a007185bc452cca227dbb215f4bc22ba",
      x"125253555245044bda38336b478b2135",
      x"af02fe1bbfd65e178495aef1acdf2cab",
      x"e409e1a6f83592efe0a0e9bde7a424a4",
      x"272da408db6f954af94ade5ee41793e9",
      x"369bc331cebda5cc16a45868497de113",
      x"c3efa04cba7dd140c1e7fafbdc1e8b8e",
      x"c9e751a6ca26f3876524a0423de00fdb",
      x"d988de06b2c89315872227d87584520b",
      x"dbaa0b3e7b49c3d0c8083c23f4c3b19f",
      x"b036e34f9f1dc42e677c3e22b91d96e7",
      x"5719802cf5c3053e782ad32fdd3aef3c"
    ),
    (
      x"f161866f029d5a0f2d8bcbb5ce22132e",
      x"a63d99dd08e8f4032857aa65304a33e4",
      x"c9260cca773f58857ba7a4481b38f055",
      x"845001960f3b47777c584be86b680595",
      x"84dcb0cde26416179b84772e59ee849c",
      x"c89dbe748a36f69db05c312880bc3018",
      x"a24cad5ad8876e5412e1d7fd254cde97",
      x"a21dad8b5e31c0f257ac0f6296a41fc8",
      x"9312dd82df89895facf88802f80bc03e",
      x"e2f874ff69da55684e38cc2dbdd28bfe",
      x"388d9e9b34fcbd20409dd4483670abe1",
      x"197cb4e987d606409c4c3d6e46de8f07",
      x"7527ff9d734d15113f8f8146cfebdf98",
      x"f4035d0da30dc988dc963b66523c951a",
      x"ace224d9b378298785d50b029e47fb09",
      x"12f9b3066410d7e19ca642f8dc401657",
      x"3b54a1fce40df4ce3edb88f9bf8c2b4f",
      x"4a09fe4ab34f1498f5a17741ec18fa35",
      x"53c29f95559cd87665b567f4e3cdb32f",
      x"2132f5037a6787b952b445a39067d17d",
      x"87961a1e795bd94a7561b641c7e2ab7a",
      x"90b348ceeee51b2ef19968945a2bb17c",
      x"ccc840ff5739411cdb357285c2e97b0b",
      x"35a29964d37c1ec6727b08f6fe178ee5",
      x"46c5381c87d3bb86808bac57d5deab99",
      x"0aa108b9a0cca5dfdeb20a7f2c486799",
      x"ea5f83fe61c7da8d0e71f05e1ceda219",
      x"2d62196563db1877bace1e649748eb8e",
      x"387aaf0ac2f5c3fd4c9fe96dbcffdc82",
      x"52d47a696515d4179cf5dfaa0e449ac7"
    ),
    (
      x"4a13d4f6a89aabdaf37c9a452865359d",
      x"1e8d3279bb8745518a25938a4cbf6121",
      x"7120a6f74eb9ac1c9c781f48a7852929",
      x"5e837e8a7a45ac5e2998e1d22c194cbc",
      x"d9265efaddd9d29b8bb87832fcd91b70",
      x"296b69ec6260e802eeef186e8c9eda46",
      x"b85ace63940acba2f4c1e4358d702559",
      x"dc20143419bc1ebd9276ab66cc26f494",
      x"59ef42d899db6746002b29342141ad39",
      x"d178cc4ca91be9c233d7835d81905281",
      x"9b562d050348f9bc4230bf6879263c1d",
      x"cc5c2d028bb262fa914146aa82e1adc5",
      x"6ae16a7f08ced85c13aff459c0840a1a",
      x"305eb0e71663409138220965ce8aa727",
      x"b19ece223ba10e7d9bad884b73de3ae0",
      x"34e0c5e1325196bc26cbe2dc07c37ff4",
      x"0f69ae903e3b1946fe4ebb4d961cc05e",
      x"01512df587a83d8730d047ba90f778ec",
      x"ee2c082ff52efbaafe8ebe5929023c90",
      x"75641a94c644f6e5bb88a5276e720491",
      x"659b90560cf58b3a2c9df533d8eb95c9",
      x"cd59e7640239951e26bf57d64b0da3a2",
      x"11c5187a64f073051ea7871d255710b3",
      x"db54c70053827f530895ec8a04a82c97",
      x"e3a69a1113d76e059be3a546ef5a7f00",
      x"0d7319850689ca80050eeebf396bf10d",
      x"b6fd4868fab069c56f378517a5eef2ac",
      x"e52ccad114782f2cbd6844c6a193bc89",
      x"1955b9851f49417538296a7d971491b1",
      x"8f9a36532f9fff959cd36f87b1b455ec"
    ),
    (
      x"3d9757c8b813f0f1c7006a389ce5ed20",
      x"9e42c255a7112b2944dce1c246d8fe8f",
      x"7e4c5b412e9090a0ab8d1f74ff595701",
      x"c4e4fcf68e94e9088f631432922afd8e",
      x"ba93f90e2eb3e0be2b30557ee89cc724",
      x"bd58f3ed2a0264a429d83398fe9b90d5",
      x"3cc9841afbb026ff0b696613b8133aed",
      x"712bd1307ae0d40805c89d8bbfab58cc",
      x"f37bc4a06dba90f3beebd7cb3e79238e",
      x"e339919ee9e7a5f7c79b60a60896b22b",
      x"032c1918cca5f3e69e1e1a9b15a7cee2",
      x"3fa740cf50c5ee7318900774ed0676a7",
      x"9c7d489183c6a1d98b0654a040337df6",
      x"20c680dbf25477820bcc405780608ca2",
      x"489dcb8c635e418ee7ce13feaba2c45b",
      x"b8e8219ec39ee4076023774a97fced51",
      x"da178bbfe0e7777a1c0b1ed0fbe2498b",
      x"ebbdc57917a240467c9ffd88d4abc360",
      x"5da20f9a960e40db5e7a2bf1e35c00cc",
      x"99df2e455fa34ac8314e5dcbdca59990",
      x"851bc4b47e4660dbf8bf4244c0e60608",
      x"4127d64091d9b0374308f0b700e96a4a",
      x"0a1380f2509b405bc3d8c290df05d628",
      x"9b09dd1ab9c1c718cec6ae18dc3cd0a0",
      x"3fd15998d6d6d95f7b5ef1ae8c29a2bf",
      x"459fff14342c1bd94770a25540929a72",
      x"5c833debe15a3f831b393f26dea67e66",
      x"b86bccd64fe040582eec8010c0de97f4",
      x"f72395b54381c3c911c26dd0830bf44b",
      x"2f251c974090cc401c2085fb5bafcb57"
    ),
    (
      x"b51176311e76848b6e73544964223d30",
      x"9963fdbb4ea7012acff856f3756b8b65",
      x"c9d1f3db4f724b5cf8495620802dbc59",
      x"8950f3796d78308a9847caf37dde7fa9",
      x"bd489106b55d1286fb1cf7e7e5841459",
      x"d46ecdd6cc0310e336c7977019b976ef",
      x"3d2e14e7750d4429a1b61714898fc2b5",
      x"b8eed0f86000f7a5c72c8fc3f03877cc",
      x"35365fbe2c37d92bfe60fa80c75d4b56",
      x"3dc48d8b2dcd12be79d07b897f106c09",
      x"f2e5144ad2303259fa13e327cc73bb56",
      x"724d53ad660c495a1291eaf1077b9f67",
      x"40b80d5be70614fdcccf84b5dede8f0f",
      x"12f9fac9a1b907fc843f4b1c080ed857",
      x"5cb89232da17f70caa111625e1b1aaaf",
      x"ca0fd233b6b9ca254cdec44fc0869ec7",
      x"a095cc9207df49b89d59a91e3a674bb1",
      x"63b37a057c7a4d05e451638032ba2ef2",
      x"4695b3c8933c05a0551fc57fa6379dc3",
      x"32fdac4a642a050b2c24d5d69b7bb06d",
      x"d1fd84226f178bf445c4c0f5038765a6",
      x"1d76b26681bbfe9a45d2644f142c3468",
      x"6795aa2e66c6b2cbd5ab42be53bc51b0",
      x"e2eef6e2abe999b81f202d577973498c",
      x"97a8cf11e7ae65bcc572e22eae88f7d4",
      x"f999d61dc6405794c3771db0ddf3987f",
      x"0328106de0bac37befc9bf890d0b0ce7",
      x"6f7a49a9c2249fbda8089afbb4db915c",
      x"fbc096dd49877ac4da028e72f884f02a",
      x"c56d5279b058cff487edcac8ac25aab8"
    ),
    (
      x"12b082142e83b3b0632813439d906e64",
      x"d59be01d04882980a48d550e772a1392",
      x"a785fb8ac1002e34826ecb01635f8df0",
      x"c54e71900371426309a2703e5ccd8a65",
      x"4d99a8e3515113113487c87d1ee0104f",
      x"e24bc0b357f3d566b7f1ae843c9d91b1",
      x"458194f50953fd6af0f0adeef6966a89",
      x"c9c78ad77763f954c30bf8aaf2ac551e",
      x"5e77a589775fc10aa06b4fb41a79c63f",
      x"4b8842dd8d5a2fe7c5b5bd91c26dd1e6",
      x"0400fc76b8ba73b2aacfd535c7c57e9e",
      x"d63b7e8049d0c5598ac94d1b062a0b0d",
      x"74d6d4135d254f8e2a1cc0d417aa49e5",
      x"6ea27f1946beebdc69953b8a3693a2ed",
      x"9c3f4ff6edaa9c492d8fb0ffd2b98d09",
      x"d37b2bdb70f2dc5863d070d1df326f7e",
      x"acf89f0cb5f531bdc6fe5d9c9aff5165",
      x"2a7bd68efc2d75d5e3322d56a2b44ee4",
      x"0931894ae15dedfb292b67cf089cd771",
      x"a5319fdb2acf40a11974b2752721d760",
      x"954f71772850ec5afd92b6e770d87fb0",
      x"07ca3019539bd63347087bd84d3be4b8",
      x"ceb2a00c0a93b476f971fbdb77ece676",
      x"f83abbafdbf79fcc22dd0ce861e472d2",
      x"e6f1f1fd7e063f1391241291087be572",
      x"500f9de6a9f681d4395214a990e1aaea",
      x"7ab041bd45dbe9fc945f8bb34c407d73",
      x"991d18a8017c4f3e6446d258affb5690",
      x"80f1d55b2e4cf3dd55cc73f836ffbf78",
      x"4eec324ce5f4fa359a3de9be0cecb7ed"
    ),
    (
      x"1b47cbf89b56bd10a67cbedd759d2d5c",
      x"4e94d35ec3a8c990705c900683423a57",
      x"1188534920e92077bf1af3ce0adfad13",
      x"85ec5a80f086064b2c38d2f8464ec263",
      x"5de53052e333a4903fd8302d580dc6c7",
      x"c7f5694719452009853792ecf70a7841",
      x"8c6a2f90d0009d3cc06ec0549b860e38",
      x"7e59606133e73221cd89df0b9c17ede8",
      x"4c1015407ac0a07518895f1028af207e",
      x"e2da04be5d7055490e8028a12752ee0c",
      x"69e6db46b9cf75a63702142c87a0499c",
      x"77c0f0807eb5faa6a998cfca5d49ff0d",
      x"280e2ce6573f76169e66558670d94989",
      x"09ed5e7c59fc35445148a374299be97b",
      x"25957e96ba130f230451ee1bdf74bae5",
      x"8bf4680dbd587d41108f7ceb87e4cb44",
      x"c6bfb5abadb84b0a3f6cd8b31623c63d",
      x"5dc2c240922fc284ae827d96b64d6028",
      x"9957ab7641caaf75d81f64eda832e34b",
      x"2e39b6e653a3aa5cb258f9210e255c51",
      x"01f87feb16f5d0c18ea09cd2a58289d5",
      x"5c2bbfc417d977c1123db7bfbc4f3d75",
      x"a3e8cb3211cf31885f268ce5057efe2f",
      x"5f2e6eed270111f64f71bcf8e2dd4ca1",
      x"25062e2685780167f5fae61f4b6d84f9",
      x"66fa01fc49741ec122701a54cf36ded1",
      x"e238f9d60e2633226a2b0ba50d8d0e1c",
      x"0d9eef26131d0824e511ed8bb39578d8",
      x"d84434b0f93794d28e85cdf31f118cb3",
      x"a8b4970a513c9219eb70cfa311586bc2"
    ),
    (
      x"94a41f0868dc485571a7c077aae2c697",
      x"344319d58d6d95a485862b31b0721eba",
      x"764a3301a3ba0719fcfd760abfbbd8b6",
      x"2301aaba85f4e687a4d0aa95e2f2763e",
      x"c0d173671124a4290d5db6a34bded929",
      x"af7ae7f57baf4c1bf4b3390e1a632df6",
      x"4aa7cc88f524bba555c3d1bff3a2a293",
      x"000410962b73fc7f810a831ab1bf0f8f",
      x"cb24c52249cdd2d81c8ca7300a5b0062",
      x"c2bedde7a57709a78cbf72ce004e60c2",
      x"1ff378ba290447c88652a3654c5f622c",
      x"365b3812c1da69b059a92eff1779621c",
      x"275ca249f6113328aca77bb3e0da3cd5",
      x"11995784e018364b47732473fc6b4476",
      x"7ca97a3bf561619ce644b0a35f83d08a",
      x"4f63076493b1a31490692ee09974687b",
      x"099e00c4bf42cb0073af685df89a826f",
      x"61d3a76ad7214cf7bacf92d33a3b16ac",
      x"13e15f3a4624bb2337f8465c8960a92a",
      x"ac1dd4f0c44ba7d5a63e57ba79a4b853",
      x"62507b26c293fd3bb692586e4b5e5fd6",
      x"861e18cb0fc67a4ad012746918a69230",
      x"a91d3e309a4ed6489edfc84ab11d8c2e",
      x"0e00d62e1082e81f17db6fc4c131fd9a",
      x"7d852490e49cc21e1e8b69a003c1b9ba",
      x"d29c8dd28eb975749f4c1c86488daeae",
      x"4eb96837b119e005c20d8b588325cf1f",
      x"f01d38cf98d22d0e2e7c1728f10c8585",
      x"849c84119b57d58a634e807aa95e669e",
      x"7c2482d38e0668426806553c373d55b0"
    ),
    (
      x"c45fbd600d2f4efa1107fdff8e196cf9",
      x"92e5a7dbe0b7f0608fe6a0d15d923a8b",
      x"11930dd65e8f8e12c706ede4110adb02",
      x"9cc914326a2e541f62aabc495278ec8b",
      x"2254242f1c3e26f92b7cf1c2e65bd574",
      x"45cea76a6ee845bfbc9af958a31b4ba4",
      x"6d731c922db52a85a70e8567a92d1bc0",
      x"f6ebb9153843af9863a4a03454df8f1f",
      x"f8b296b72d01d9fb6f38f62a7c5fe3b4",
      x"3cacf11ef295f028cdbec5771ce1c04a",
      x"d0992eee4ec698a7013b0e4723f508f2",
      x"32e37b0275b533da061cef54c8a1a767",
      x"1678081a1bd1b0c00d8010743d4edbaa",
      x"bd0fd8a1bf354cca158bd417d8ba5bcb",
      x"3048dc9c95d3b37be4ef84ba716e930f",
      x"3f4b99cc59193432192f035b12f6774e",
      x"d8e34ba397a9cf7250bf0481c5a80cfc",
      x"fc240133068ebeb92957399b78466f58",
      x"06d5e595c921736f1b1ad83af8fe203e",
      x"b6a536ca2a67ba46f67d656df909a543",
      x"9bf35bc3999cb49e73a590aff9df334e",
      x"b0dc980c6e6146a181da04f557d76c95",
      x"b8a2af5de9341ac4663264fced54ffed",
      x"5cc35884288e5024239ff03b888b93c9",
      x"6a9ff1bb0708de3261a1f9199653f204",
      x"b3dc5123bdec7686829eb072d9a321e9",
      x"1c3d49fee69a5ef53164e4bee1fef1f0",
      x"b8364a8d97758423a39841d9c5efcf1e",
      x"4b59daeae8af91a7a925a6d2f3f3c852",
      x"25bc7c8d680044f137d8c121c7596981"
    ),
    (
      x"2dd10107f97e5de6afda681f7a8ef49a",
      x"d337aec3c5ea7bb96ef1fa61d0c6ade1",
      x"698b24fc15daeea4e9f6615b6bc54dc0",
      x"6a4a93bee6eb3e9595284c337692d4cb",
      x"0213896a8831e72277b744130f936686",
      x"280a58080db0bfdf8ad0c7408973e872",
      x"9ef214bc8926acb24ca87cde73f37e69",
      x"b91f4debf8ec6c5e53c2f84919328a0d",
      x"a6358974664262a1b432f55c299ecfbd",
      x"4b587c3e3bb7f9ecfec0095a85110e5d",
      x"59cda7bdef604b481b13003a74890153",
      x"ffc0006584680a85c9e63e62857b32e1",
      x"f5f957f8cd8d26995789214ea028cadf",
      x"9c018121b135c6a9fc6e096cdcfe875a",
      x"da9d867c0f6c0d32a3eeeac8fd95991d",
      x"bedaf2dd4d4b934f19ce8c083d6c5288",
      x"41b13298ba4ded1f6ac6f38e5fcb51e7",
      x"92032d218bf3bac7c4c0d87e01a2b4c4",
      x"4fafe0d8acfda09b6085550a817e279e",
      x"c0a7c95df5dcba2193a223353d4e6b61",
      x"67ac9c8a0f4f776a21cd20f69c8bb84a",
      x"ebc226ddb399581f9c432a0db378ebe8",
      x"11c82e55f89b550118864586fce6ae32",
      x"a7e1c8741588a77ec2b4b385b065cbfb",
      x"f1e57159c0a15bc67186e2fe41dfb48a",
      x"f74dd81a85fae06ddcb91dbad9097d27",
      x"a240a91812efbb6511b7cda979e7da02",
      x"811cfefaa031f7676618455e1df2aa54",
      x"9ff4d38294eed41ef3502793b4849074",
      x"76e899b12fda1c75bc5232f8dbf48dbc"
    ),
    (
      x"7b999412b7519917fbb06fbad7be157e",
      x"a509de8d39c603267e12a8bb528be74a",
      x"9da7a74a476b95c65f10779fa12493cc",
      x"0e13d0c8f97b1bf07d9c6d70356110b4",
      x"b1dcef19ccafdc806bae7e7d731744ba",
      x"6ce582c7b30adc05cadf14981526cc8b",
      x"a08ca3033a5fb2f11258ca3ee7d2f2a6",
      x"ed5332e3c9f43dcb1d74b2ef1045650f",
      x"0537a6d6eda2452a61249fe3db98028f",
      x"791c7d1f1952b3337a6dea5b3978b1e9",
      x"f79593f3b76dbddf1d0ff34885d19ef8",
      x"ca87906815059248e07b36273f50217d",
      x"f104814c0d0c315a1fcecd669c12188e",
      x"cc455a0a9005e388605a8aea7fcdc73d",
      x"5dfac939bfc2c597608e714a79de8e4a",
      x"3209fb07044b44087be2a4db925c83a4",
      x"7c04080b8badb2f0f11876f1abfece5f",
      x"fb92d2af29876ee79ceca4e8f7d103b3",
      x"ea86f627b0798cdc3f46963b74a72990",
      x"7522b456dcf5e72e0c60ec7420a29057",
      x"477eb6e2e5f2d65839b4df3030afe3e0",
      x"a7ddd0272a6ed96538646a562afed3dd",
      x"d61b25b698cc04af4cdee78fdfc7bf3b",
      x"0b0e54a0ddfdfdf1cc472f6441175665",
      x"986ca56a1a8a23d879930821f54d7110",
      x"64211eaf8f7cb28efef53ece1fb19966",
      x"9534818ce58ba6238f60dc2dcce19c85",
      x"63b34eb48a4a4647d67fa2b384c48465",
      x"ec4b357bc64e03497b3cccf6f5f56cb6",
      x"edc136ac42cb5d7fc079558c8fb6f940"
    ),
    (
      x"5e8bd598592782394aaabf1714f0c896",
      x"aeafe5efa672efa6ffc2051f4b56e261",
      x"2ddf566d5050c72cf29f350644c62e9d",
      x"872343789554cd5f2857838c1b6882b3",
      x"2a141672f58722c102df11ef1dd8b9e1",
      x"525d3783adea2e213c5e2ad26e43123f",
      x"b952db9c5169de42f1ca7d8b9c126b97",
      x"07b7bc47ab9a5a2b4f6c8c87161122f3",
      x"e82531bd0e5d29dfbbf03d1794d7accf",
      x"10135abff2ca989ee81de2343a5d9098",
      x"83a4dac49ee6567c38709c2ff840a910",
      x"edc25c4a3a9cbe3eed878a693314fd89",
      x"ed76d9d53342f1abaad06fc4032b58c8",
      x"dafb50ce9e890c10dbe00070d32842ce",
      x"fb2f0d5bc2997802afac4352855dfdce",
      x"217fcfe69238f285fe4342ef1ecf4c0e",
      x"6cfa377fff603695d53eb77620c550ab",
      x"e0722272d54e30cb1f62a51f88377a53",
      x"0b13cbf5087af3a5a1ef0dc9389f9f31",
      x"69a8ac4f8b1e788a57e6fc7480a44086",
      x"be7865566bafa5b1b4b2000eacd00f0c",
      x"5c86b22f6cb7ec286238807e91a3f925",
      x"e1c8f7a190d45c2a1bb208f03606162e",
      x"25312b407a27413d026b5966901f0908",
      x"41ae15e146d679a7406c43dcc35fb2ac",
      x"f83dc4eb84e04efb28e9d97f66c25f4a",
      x"61d83644e4988007ab71abad818907ab",
      x"719bd08984cdbac7058f3e7af2ca1fe7",
      x"6da878c0ad93ec5768f40e906f5a1992",
      x"50783247c565e1bb80c6265da3d19210"
    ),
    (
      x"43c602b483ab61e25af0b15d2fe5b6e9",
      x"505318798ee0216d44054097f11c9ab0",
      x"11ac5a3e3cc1d002a21fabf5d3c181ee",
      x"4c7cf9737d643ebcc318d1460182d5cb",
      x"4c2415a7add26b6103bc3301e9528290",
      x"c053875d7e91a86378f2d3557e68ec25",
      x"b0987cbec0c7f820fe207592b1438fe2",
      x"092ebab241eb53817ba88ef8d19e8d95",
      x"6ef60fff7ef74d62040b0149a8720b78",
      x"0ccdd6969b9d4c65f0986a8cc3ddc157",
      x"072de58191d311bd0e72efc4b2b1fdbf",
      x"99f5114890ecf8619ffcb861e2f895a5",
      x"f667cb81af391eb4cfc0a6a43c5b6565",
      x"43b71b40b2f229378cd1df9941ca7b2a",
      x"243f630201926629dffcf1c8edbc4337",
      x"272c086cc836b057bac64cb4d61e67d1",
      x"5efe619cb2faaf4513c3cef6bb67094b",
      x"f5021b0425915b1f22d6019debcf892f",
      x"649ebae5474d7e85ddaff312f303fd1b",
      x"18627bcde5e5d2a0dcfb1778f4820803",
      x"133bca4374722068cee59731ecba4d16",
      x"d70ed0c4e186cc9ab006732f04bedc0a",
      x"cab859041a1e8106bc373ae6600c479b",
      x"ecf101ce2ff3f7074577cd7b2045f4d6",
      x"c52cf9fd9f6c9967daf4d026cd9753ed",
      x"4399792dc6aed194716c5ce52303aa25",
      x"2401a10f98e0d19424a150f16380dc81",
      x"c56811b663bfd624bad79918211f81a7",
      x"610081f27d46bbdbdff2b7aee63d8cb3",
      x"b1f2cdf93623448fae0586c24d5fd8fa"
    ),
    (
      x"a192a8db4be2bf60d579a5ab910e60ff",
      x"70aaa7d5600b4e35f249d480bd277a35",
      x"5bab77cd83e6aef25ed49e949bbbd3c2",
      x"c77fba612cbf92322bbb18909c0db96d",
      x"3114965eaff8ca8c548f31109f346418",
      x"a462b94b466f2406d6cb02d3374ad16b",
      x"f86d18b50a2980f75d97a54ab8113f04",
      x"9078c09f9fca82cb4fe1d6d2b2921f05",
      x"f5aa44b13859e7ca3d599bbab30c391a",
      x"6635ae2dbeeb3d971c280f5b98b2bdcc",
      x"9875dc6f85b371df01bf4402b2bb8c12",
      x"25bbbf8247d27f57e23602240689b44f",
      x"4b2e1541c6a3536ac03192047a3dea54",
      x"2ad453b85206bfe17de6d7c37bf2af00",
      x"bef894849e67f2c8f988647fa07dae5c",
      x"09e4b3dd016d83ca208627bf1e5d1cd4",
      x"7a26d6f90e203f36c18f27602d3a4c3c",
      x"ae394e3cf0eb3c1435e60418253d2900",
      x"9c6f42af4448741043a91a9ee89323a4",
      x"5402ea88db6671eff43d33d33939a1af",
      x"5c05a9717e347b725e7ebcd3d58498f7",
      x"63cae68264dc07c1c256dd1aeac0e983",
      x"1017228e6448ac19c39cdbe6a95c6472",
      x"b7bcb333ff22cf149d971a3909e18842",
      x"497de27408a22122c878fbfae185239a",
      x"5919c0b9195b0d88e2fb8bd81bf26f24",
      x"d173411f0cec7c3b318fe2e7538a7900",
      x"ad1e1b56d19f52c0bcee477b2a0df886",
      x"05af863d9e1de6fe166e343504a48f21",
      x"e5a016f041630954cb6a5f409178e85e"
    ),
    (
      x"5e2e1c72bb6942104c74da4f590cb8cb",
      x"3b117160a8724a8a644c03e5b73090bf",
      x"e4aa2dd4a740083303ba1227ee3d3c9d",
      x"3eee184a2a1e072b099956880ed894fb",
      x"a8f5e63ef4526212363d02e4feaaa3ca",
      x"bac342226779d19434a7d271a735fea5",
      x"04c55f4edd7917de6151070f7eabb7fb",
      x"c046cba1d1dceef743c0ff7d9fbf5b58",
      x"25b426735becd74efaaaa88a42092e64",
      x"1fa995b4d4bc6601b1236271d1103d7e",
      x"c2e42e73bb2df12812bd8039ab054485",
      x"00fdd335d2e4dfbbb1cbc6f39acd2e65",
      x"2f32a8cc5860d3162ee2c33b3fc23774",
      x"b1ba18342fc78e28ffee1cb468dbf524",
      x"b8b9d6621e227903ce7473ffa6d0e33d",
      x"a0ac4e5a321439b944f508838f736e2c",
      x"6a174bcfd52ae40f36fa28ed6462be70",
      x"7a2f0493bbf396c6f24010cbf55551e5",
      x"65171b3b5980ba12c31e055ffd8340a3",
      x"b83ac3c41b82fa45ab9d84f5c141840b",
      x"cd602d191e8d389a0a65ee0a3cfca630",
      x"b1537bf46606b0a5f85d55add34071c2",
      x"c6919b90f5dc26f4183a91eab3dd126e",
      x"6c24a4aedff7ef743ca473365701ffce",
      x"1ac7707368962b0d38d90a610058d1ee",
      x"76c25e92f66be0237ae5cfe623b5b406",
      x"7ae1e1e1f77608c447ccfb30cfde68f6",
      x"c302fbc872fcc7fca233d2fdf231214d",
      x"7e26dc1a2cd05bca66a5a8e07e3d9ea7",
      x"7feeaf5f9011a66795dfb3286e2589d8"
    ),
    (
      x"33a0501b6b8b9767d6145fc2be7ea651",
      x"c846799c838e48373cd6d15793c7b374",
      x"23b68b9941228749da9124870cd8979b",
      x"1a4a26564fe1762907015ba7c7e83c01",
      x"560483bfe1d5aeedc9a85fbc81663982",
      x"5dbf12af3114e7074066f91ffff3eb05",
      x"f10d01418fe75bdf4596adf7fa536290",
      x"0d1538efd7d51383009cfc615e2872d8",
      x"2bc93ce124d0e237d546210be70a4376",
      x"f27834b7869bb382e36b5a1bf9c9df2c",
      x"863f3521c107a91209f5999e11845395",
      x"384b9ed1a5f1df9525e18808fa7b55ba",
      x"3f49b821a7582bf258cc75c50802d332",
      x"fa3fbff509fd1a806a7d45dae9ac0d12",
      x"8198d91d3095a562b28c8465ef77cdfa",
      x"634f84ea6880dec7205b30aaadda248a",
      x"a5ad7996932a54f724f4d98719ab3f0e",
      x"bc17483a1a549ad024a0a4375ffa4e80",
      x"48210034ea736061c232e7729dc8898b",
      x"cfaf3b6d15cb30f7a15bdc9a2f6344fd",
      x"319382bdc8f81d04ecc79fa56e1c7609",
      x"a63d455125002149534240be776a43a7",
      x"759a2e5f2bbc6ae0dfda08906de31266",
      x"30389539e00d5d31c847cb86b3c786b6",
      x"31df182c0f548a111ca8afbd083f3888",
      x"363702a0c1b0bc2c01963328581f1c1e",
      x"8a752de050d83b4ad1c5b7ca50cab929",
      x"a8b7e8f862a9ad63bc2aacc8ed6a85d3",
      x"00a3f928dc69210176b9b23565abc255",
      x"caec1394f20dc5b8b594bd2ac9a2311d"
    ),
    (
      x"2c16e35160299d76c19ca7fb219f634b",
      x"79fa54af2f38e0dbc48f15696b7be999",
      x"8b9d422bed2d8d84941579b38aa491fa",
      x"bcc38b2f4db13d776f6bda9adebf217c",
      x"34238118d612603bd56550b0bd267350",
      x"cc542d08860534c239102eda437b6768",
      x"feb789e3e1776ed2bc4b337b073c4748",
      x"bdc1b7bd990f482a849b67fc59dfcf5e",
      x"ca01b071e8c8115af01331969f6c4394",
      x"9148d3658d5cb00b8898480cd8bf47dd",
      x"690ea9f82e6e183d1c162e37db3d3b99",
      x"15fc85c4d66ca4c6607000eac4424de7",
      x"8cbe35fef69c2b04e131a65eeaed005d",
      x"213f0360318d844475507c106b813397",
      x"dc203c8a6429dd5c6bc2920d3a241c9e",
      x"a6b4bb569499cd06dc26f5b46e55b17a",
      x"78ef3101d4f019c866589a4d4abc688a",
      x"d1ec6e7ad39a0f7f73d0ee19b2771d33",
      x"531112577cfcc155a91de7012901ef9b",
      x"6fa7f78a272ff33f9e2f47547c4646d6",
      x"990d5fbded30dad47938d3b58b57d9d8",
      x"718a919839d0afe7875861c0d269ba0b",
      x"1aa139b72b08ecca5fa889d5e071eb8e",
      x"060330e6b4b82d3802aba5d9de27764e",
      x"92b325cdc8bf69a217fa79a18eec9973",
      x"3572db71046922453c55f8740413e595",
      x"cb319be40cb892278bf80095b4908c08",
      x"4a1113623b428166d8cea4549333b381",
      x"adc3183f0dbed6c9519ce796f3a29891",
      x"1bf3f9dfbe0fb04c16f14204b2ee6bd9"
    ),
    (
      x"58fc3107b6bbbcc18fb46551086c402f",
      x"d7a41751128fa928563e06b3dabe793e",
      x"82ef7ef9d5e6c0245867c01cca276b07",
      x"08edc759ff1d82f31a2815bf5fb45bb4",
      x"e4a300e3f82b9e414cdd9bdec36e7002",
      x"a37b50a6bf55a19d88531ffeb186c6f1",
      x"b905804cb7485874e0578c19883a4cf4",
      x"0bc4b6c12f4d4410b3335e59dc35d38c",
      x"13c5d7ac8d591fb9049c1b31574b82e9",
      x"4635faf51dd6e6c214b012fa831ffafa",
      x"30e3142f8eedda1de8bb51b493db1213",
      x"b2bc420f7857f0b77a58d5c5f9fb0d55",
      x"5aa19bd7ef13a10b036d8ecc4bf5cb00",
      x"a875794c6fa0990fdf5e96efc76e8b12",
      x"5c2c5ec90797722412c8302133dab0be",
      x"290680c83c0cf88b9c7f41b586ca5be7",
      x"5ed42461b85f093c2cfad3fc1f1cb8b0",
      x"19de7cf2beef6b6ef24a5c11b17db94a",
      x"cc60f5440d2b2b637356128b35b5f8a8",
      x"b5d156a1f1337b1e27a9c0678e57f032",
      x"70d77cde169f684137914bdc9f6262df",
      x"0d4aad73531ba04683accc449fab78c0",
      x"c03c6531b3e62cf1cc31a83bfeb45e74",
      x"0f45c22c556f1f21e6ff3b841a68f9bc",
      x"65b1f37f1c7ae00a9bd4d0f38e9eb7ff",
      x"68d86c9a416ad1b03c9f0f2d5cada782",
      x"52b188e99632920a2890784a31efc409",
      x"e40e1fbd94827b0a785db1e58f74cb99",
      x"85c9d5be685f9ae5a7be3083fd7ca936",
      x"5101e09abb45864ab433aa3910948e17"
    ),
    (
      x"a3872b92d9f16ca4be968fa6b9eaeb29",
      x"d986b4777c7ece75ef1e63f767c537b0",
      x"a0468ef6d6c54a4e5ba966c086714c63",
      x"268c7700f77ce89371ee5400ac54ec95",
      x"84290d421796e2c042b11c2c89c85535",
      x"c7799cb53d2409af3ced979ba78f7da5",
      x"308f6df52c5b602c45986e4d689d379a",
      x"c0a0d8cde7d0d9d6de895328d91270a9",
      x"8a878a0ec9a4bf13bc00870268ea8298",
      x"957a58b307f36a006ddcf599c1cfce8c",
      x"e885a5bbdfccbc592d7cc5f1741d4097",
      x"02e19083db8bd854759de79247472613",
      x"77566ad483833d99a7a856d0109e42ed",
      x"eb521dd6cc8725586d94376094becca0",
      x"f1d6026a253016bde66b99fdb19d1953",
      x"6beb6b0ced02436d16268d010cfb3bb6",
      x"50b60b37b9e8e9983aa0177bc0fad96b",
      x"f55daf22b96c8d658d37b1bf03cda5bb",
      x"80083c2cbfdb8241d4f1af1ce07fe768",
      x"61b07bf1135442cd403ddbbf93106510",
      x"dfe662163b52e99489e5c48c1b55dbd4",
      x"d27f78fffabd53cf2989b4abc62d2973",
      x"e69f22fa3cc8e39de19ea7d01a9ff1f4",
      x"352de037c257d17626b33b168eb318bd",
      x"5d6670b73ed97ff3642fb68170812db3",
      x"91ebe4a0df0fad0bf536edea9f87e73b",
      x"e029149a1cc91a37e20c64fe4d350d8a",
      x"5f361792807912bd64885f9c0fee6455",
      x"b7e9ec0fb8228256dfe9f6add2a79004",
      x"cd6d900fb99745dd6f25231fd9cfa76a"
    )
  );

  constant ZR : T_NN_MATRIX := (
      x"a578bc2b1ddc014f9cd9591d22768177",
      x"10ab610fbad4ce0951518bed0f94a067",
      x"472021754963d954918327fae562262d",
      x"593628d254ad954c31dc06ce14da2f3d",
      x"add61494c765a0a06c5802090f067635",
      x"7d9f9925d602a1b76e56850dc85da44f",
      x"8aceb851ffcf77e4e86d91f7cd530af6",
      x"829f47a97839fabe9f3fd90631b0ff10",
      x"0598fc8af0f8219b08b89fc3efb9229f",
      x"a0c57ecb8d33c99611a1b26fd927d774",
      x"4f695e0d730050674b228f123a4a257a",
      x"ec1f9e6ba954217c0993b047a0a3195c",
      x"1dec62ddabe3f0251eac2d3f201cec7c",
      x"330f427458e8c989eb7a35954b201f9b",
      x"4130592606cf19c2e0a7cd47bdf4ac84",
      x"6f17d5863f332af48e94b02f66bcfa13",
      x"46f9e496e175308c7512f04fdcd8ae45",
      x"9ff3491612ed9b2766cac62b9159c0bb",
      x"5aee5ef2c6ba96fdb6bc94b241b43fd4",
      x"d1b15866a8324637d9edf62e8ff2ac36",
      x"f6971ee78b44fcc4db2251548b499fe2",
      x"7f959607eff2dd0bc342a99b552a6ba0",
      x"a6b29630a7204f545432d83e4899c809",
      x"b527a180d561ea0c9c7956e878c8f7b7",
      x"8fdc55b2c60d24e14a138b6489b929d5",
      x"2078ce8833849aa7fe308fca4299a37c",
      x"22a1a3e43fb7b55febe48b5d203e8fc3",
      x"227e4e8ce1b7ed88d4fe7afdea4f0e55",
      x"d30660fdec3896b959547aaa1071c2bb",
      x"a7b48af3be5450e6bd9d2b8ed7947be3",
      x"ec94db899a4326ffd0bd7a2f50f17429",
      x"1f368a526f1b10b3887f6a9e8b68086e",
      x"328cec75dadceac260cc474c02a33d0e",
      x"d5dcf224845d00fcdd58b5aa17e32ed1",
      x"de3e44eefae105c272f3f948c571d0f7",
      x"55ec9e6ebbfdbd85052375438a4f3a21",
      x"f384012ad3407832e27515b8f6d7d9e1",
      x"5e090ccf7bc12792fe4fe2cdc95ab1b4",
      x"afa5d9bfdcbde35c7297d08522aec290",
      x"c099c5175f70807e3e0665812513bb79",
      x"e62ef51f278b17b17c463a5ccc20617c",
      x"3ee1a3ed71d5d5c40f0dc73e531dd175",
      x"b9b094bddd0b32d32e04a4a6af488f87",
      x"b82aec9038924ad86eee9419cb1b4458",
      x"4297c5059f054b8cbceb1eb639ac87c2",
      x"1e9696f8ac90ed3ab6e5b8129cb1fe94",
      x"81db8c6aef67e46c12af916413f163ea",
      x"4be92507935db35257e3c2ebc307422b",
      x"fba26eb970a2f69389481c13b6302c49",
      x"d053e5aad8df4472c5afda53a3282716",
      x"cbe000839213365e69205075b270dfa2",
      x"4d8a51b67bd4176e53a01119368a878c",
      x"7e41c4ed8001abc8582ede61956aab48",
      x"61b363c6ee0568eedb0859b7c9c0ef2d",
      x"ff9baf368782d726934ec3bea0bb93c1",
      x"4bfb1cc6aaf85b4d195d62dc52933d01",
      x"999705fed878ca1c9dfa476d854b1453",
      x"4fede96508963e0f95fcba27779ed84a",
      x"1714975acae8177b5a9579ed7e997be7",
      x"ae2fe46d9ca83be4a6199650979c0c41",
      x"d7d024ae61c86e699775b974d7e673da",
      x"a0df04fe5986cde5d15801debd205413",
      x"750638699cdb84207834ec8f4681414e",
      x"083fff970d6f7c8138f762f6ce334b62",
      x"9a35fc2a6fff039855bd01df0b49bb13",
      x"44b6eff1fc5922e98afeaf2bc8c8fc25",
      x"0b08e62ca8460a3383d48591c409e810",
      x"4afa713626a3fdcfeaa9e803d25941aa",
      x"92503ee6216ac27bb6a9bdb82c3a133d",
      x"3075649fdb0d2ffdf60891ad5d2fb84a",
      x"a35c8896bcd605e2c40434f5232ea82d",
      x"98a67870d2bc4f1c8a6481eba1d45e21",
      x"771e1fb20e50082752a11e23d99369c3",
      x"5b2debf63ebdaedf28cc0f676b25a233",
      x"fb907d83b372b2640d0a439cf275ed04",
      x"b59ad77a94d6e43fa02c7be7fbc07166",
      x"6263b3dcc2ab6ff9e8feef8a137e43d2",
      x"fd31be7b78126b45c94fa78a82de7780",
      x"648500fb6f12204de1f14d6220d89cda",
      x"d9d32f9c506aff987b6eb8de1124c997",
      x"076de08d0b026af00a4efff01b2eaca4",
      x"cabdb1d7e3f788453c5823db3df8df30",
      x"986eeedee62a47509384adb0c5da9bcb",
      x"5aae7c24f2766a7c408a8c8d623d1160",
      x"d5db86a650e90f32b356c5b3e738655c",
      x"fb478b4c7b8ad32bc57c66cbaf4b31ec",
      x"a4f19014023d51c8a3bcf10f095ee6c4",
      x"2928bb2acf89aef0628fda27c18c5731",
      x"61287e76d1a6e9db28889ee31e545b10",
      x"e35abc245f7a023643e76b8e7aabceb2",
      x"e094a7367b60f6317c86aedf8b8925ad",
      x"99848ddf3121c2954c4c0d141f48d308",
      x"f0a4409736f625b65c93da169f79cb34",
      x"9f5e2e1825e2101695d121fb3608acb0",
      x"23792cff52022ac96ad914154ea6e620",
      x"b7f1b8f871708b88b7b861cecb2af39d",
      x"8e5a5164cc3de0ec619765db85d5f942",
      x"1fee498b53ee63862d4b3533ec136941",
      x"6c8b9dc17f1e6ead0def8258007de0df",
      x"9efa17f4e1335bbe0bee1ccbdc6dd9d0",
      x"2bae1ab09b957e453182160e3bb562df",
      x"f897dadffbd737c23f9b0924556744fd",
      x"5f741e6ec74e7d5acc9a5a2b621a8d66",
      x"68fa3ab9cb83b46a801eccca2de66a22",
      x"0f71ea99f7265ede719d4c3ecc4503fe",
      x"2de5812a4b7a29eba35288ed7468e2a2",
      x"afbd53d89a1cfd1d78779c1d7f627e2b",
      x"c3c5a6ef4d55eb382dabfe763c85a6a1",
      x"f045d31888fff0535b055fe76e7ebff8",
      x"234bdb9dc8ed90a26529bf9092a76d1d",
      x"c0bd1f2775f8ff5363910e13cebc6da9",
      x"a7c9bfe618bf83794dce5ed72fd2c55e",
      x"835d902cdc3dfc4603521a5b926afad2",
      x"696bc7ea5636a30b1026311fb955c9e0",
      x"c56f03b9c50992e3b9e1a4489ff2f7c2",
      x"556f49d077f33f922d2a12ffa8ecc272",
      x"2c5adbd7bfc551534b84f8e2950ce61f",
      x"4abe17140e16d52637da1e3e8d6f2398",
      x"d55af7e8596b51eb874ab318dc27255b",
      x"67d2c514f54874f03d4d4feec31db827",
      x"bd376e95301bdd11304b7d54224813e4",
      x"de668873e4bcd7707d62f064a2c3b869",
      x"9a5dc3dbabe9a62c5e3f584da0009322",
      x"f38ccaf41bff9df9b14f87555c18748c",
      x"27eee3bc8baae6dd18b650489689b688",
      x"e983f71844c053f199ec52153654b371",
      x"80d7a07887b61b9f856f27fa16f585a1",
      x"6c59c7487e39fa98bd07f4a5906cfbc1"
  );

  constant RMATRIX : T_RMATRIX := (
    (
      "110100000010001000101011100110",
      "010010100010101101111110111110",
      "000011100000101111101010000011",
      "110111011101110001010011010111",
      "100000010011110000001010110010",
      "010001111000110110011000110001",
      "101111101110000010000010011100",
      "000110001101110100101001101111",
      "111101011001010001001111100110",
      "001101011001011001011100001101",
      "011101011000011111000101101011",
      "101101110101000001101100100010",
      "000110010001011011110000000110",
      "000100110111111110011010010100",
      "001000011000111000100001110101",
      "001011001101001010110110101000",
      "001010010111010010000001000101",
      "111010001001010001110010111011",
      "001100010101000110100001101010",
      "101011100000010001110010001111",
      "001100000001011001100101111011",
      "010011011100101110001001010101",
      "100111011011001011010010010000",
      "011100110010100010000001001101",
      "101101100010011000111000100101",
      "111010000101111100010001011110",
      "111001011010101111001010011110",
      "001011001110100101100100000111",
      "000110010111100011011101001001",
      "000101000100100100100100111111",
      "100011011000010110101100110010",
      "010110110100110011110001001110",
      "011100011001001010111000101111",
      "010000001101010111011000101100",
      "101011111111010001010011001010",
      "001000100000111000110111100000",
      "100000000110110111000001111111",
      "001100101010110100001011101101",
      "110000011110101110000111100001",
      "101000111111000010001111111111",
      "100000000110110010101101001100",
      "110101010111011110111000001111",
      "010100111111000111100001010111",
      "110000011000000010011001111100",
      "011101100010000001001001110101",
      "110100111100100011100100000110",
      "111000100011100011010001011110",
      "111011101011100111011000000111",
      "001101011000111010110111111010",
      "101111011101111000010100111010",
      "001111100011000100100101010000",
      "111011101011100110010110110011",
      "001001100010101001000100011110",
      "100100011000000011110000111101",
      "110000110110010001000101101010",
      "010011111001111110011111110000",
      "010110001100000111010010001101",
      "111001001001010111010100000111",
      "001011100010000011111011101011",
      "000110001111100000011011011011",
      "101011001000010110001111110100",
      "100010000110010010100011000010",
      "001100111001101000101000000111",
      "010100011101101010101010000100",
      "001001100111101010100101000010",
      "110000111100110001011000000111",
      "111000001001000010011011101100",
      "100100101010011000001000010001",
      "101111000000011100010111000101",
      "100101101011000111111001000110",
      "001101000011101000001110100110",
      "101000110011111010110000100010",
      "100101110000000110000101111110",
      "000000000110100001111100111010",
      "101011000101001101111000111001",
      "100011110101011001011011010100",
      "011010000000000001101100010101",
      "000100110111011101110111001101",
      "110111000010110011100110001110",
      "110010100111010010110110011101",
      "001000111110010100111111111110",
      "100111000010000010010110011110",
      "101111011010010000011001011001",
      "010111100010111010001111000011",
      "110000011110010010001000100000",
      "010101010010000101000000111100",
      "100100100110101100001000100010",
      "001101001010010110100011100101",
      "100111111000000111110000100011",
      "101110101110100100100011001111",
      "000011101101001000100100001010",
      "111110101001101000010110110001",
      "101100111001010100101000100000",
      "100110111111011010111000110011",
      "000011000010001100101101010100",
      "011101000101001001000000011100",
      "000010011111010011110000100000",
      "110000110101110101101000110000"
    ),
    (
      "011001101111011110110110010011",
      "101100101111011000101101111011",
      "001000001100100000011000001110",
      "000101110111001010010010100111",
      "110100101001101001101100101101",
      "010001110011111110000000010001",
      "011110001100100110101101001000",
      "010000011111101111101101101000",
      "111101101101110100011010001010",
      "101010111100010110000010011011",
      "101011010110110111011110010011",
      "111010111110101001110110000011",
      "111000010110111101011110110100",
      "000000000010011000011001101011",
      "001011010011011100100000110110",
      "101111000101100000001110010101",
      "111100000111010110110001011111",
      "111010101001000110001110011010",
      "010100011100000111100100010010",
      "101010110000111110110001111101",
      "111100000110001111100101110000",
      "110101011000001001101001101000",
      "001001101010000001001101000111",
      "100100110101001100111010010101",
      "000111111010001101001110010101",
      "101110100100011000101010110011",
      "110000000110001110111000100111",
      "011011110110110011011010010010",
      "011001110001010010110111110011",
      "000001111000011010110011011100",
      "110110101100110110011101101101",
      "010111010110000010110101111000",
      "001111101001101010110001000101",
      "001010100011010001000000011010",
      "101000000111101000011001110100",
      "000110001110000100011000111001",
      "010010001001010100001011111110",
      "000101000010000000111011100010",
      "011010100000001000110011100010",
      "000011001000011010110011001101",
      "000001101001100101001110010001",
      "111111010000100101110000011011",
      "011001110010011100110011110110",
      "101110101110000000100111110100",
      "000111110001011111100011000001",
      "011011011111010010011010010110",
      "101000110011010000101111001101",
      "000011110011011011111100100101",
      "010101001111000010010100010101",
      "100010001111110011010001111101",
      "110001011101111110111110111001",
      "100111110101001111111010101101",
      "111101001111000000001110101101",
      "111000110010100010001100010011",
      "100011111100101110010011101110",
      "010101111110011100000101111101",
      "011101000010100010111100010111",
      "111001000100111010100101001100",
      "011111001010001011010001010001",
      "101010101000111111111010101000",
      "101010110010001100100010101001",
      "001110001000001010010010000011",
      "101000010001011010010011010000",
      "110110100001111100010111000010",
      "101010010110101101001011101001",
      "111100111101010011110110000111",
      "100001101010110111100011101110",
      "100000110111010000100000100110",
      "001000011101001000010001101001",
      "101000110111111001011000110011",
      "001011010110101110110000100011",
      "101000101100010011001100111100",
      "100111101110111001100001111101",
      "100000100101000110000110110000",
      "011100000101011101001010101011",
      "110110100101110110101001000100",
      "111001010001111111011110111011",
      "010100011001101000100011011110",
      "011001011110100111110001111101",
      "111111010101000001100000001110",
      "000010101111101101000010110000",
      "111000001000111010011111101101",
      "110110101100111010011111100010",
      "101001101100000000111101010000",
      "000101110101101010100000101101",
      "100001001011101000111100100000",
      "000001011110001000110100000000",
      "001000100100000111111101110110",
      "000001100001011101010111001000",
      "111010101000101010010111111000",
      "000100001000101111000110100101",
      "111111100000000011101000011011",
      "111001000100111010110111110101",
      "000000011111111100101010001010",
      "111111100001100111100000101111",
      "001111100110011111011101001000",
      "110111000000010000001010001000",
      "111101000011001011010010100000"
    ),
    (
      "100111101111100001111100110001",
      "100111000000111111011001101001",
      "000110101010000001101001101011",
      "110001000011011101110100101111",
      "100000101011101010010010101011",
      "111001101100100101111111000011",
      "100010100001110100110000011011",
      "001110000011110111011011000111",
      "001011011000110100011001100101",
      "110101000101110111111000101111",
      "010010011011010111000010100000",
      "111011001001011100001101011111",
      "011100011100110000101101111010",
      "010100101010010110010000101110",
      "011100010101001000111101110010",
      "001010010000101110010101101010",
      "000101101010100110101110111110",
      "010010011101011100101101000000",
      "101101101000101010101101100011",
      "111010011001000011000001100100",
      "001010011110001101101001110100",
      "001011110100101010111000000110",
      "100010101101011001110000101111",
      "001000111101101110100010101011",
      "100111101100110001101111111100",
      "110110100001111110000111000111",
      "101001110010001100001010100001",
      "001101100111011110011001001101",
      "100101010001000111101110000000",
      "000101101111100101111001110110",
      "011100000101000100110111001000",
      "111000101111001001110111001100",
      "011010011101100001110001101010",
      "101110000111110111000011101110",
      "101100110010011111010001010110",
      "011001100110111100111000010000",
      "010100000001000100010011000000",
      "011110101111011111001100011000",
      "010001111000001111101001010101",
      "011000111101010011001111110100",
      "100110000001010000101001101000",
      "110100111101010111011110011111",
      "000000110111100000111111100101",
      "101100010111111101011001100101",
      "011101010011010111110110010011",
      "110100110110110111000000100001",
      "011110110001110000100100011101",
      "111110011101100100010100101111",
      "110100010110110010111000101100",
      "101111111100110011111111011111",
      "000110111111100001000010011000",
      "011010000001011000000110001101",
      "000010001000100001010010101010",
      "111100111101101110010001000101",
      "000001001000100110100100111010",
      "110011000111001110101010110010",
      "111001001110011110000010110110",
      "100101000010011110001010100011",
      "001011101100111001111000011111",
      "101111110011001011001001110110",
      "111111010000001111001111101011",
      "000000110000110001011001000111",
      "011101101110100111001011110100",
      "101010111101100111100111010011",
      "111010110001101100010010111101",
      "001101011011000100100011011110",
      "000010000000110011001111101111",
      "100011111100011000000101101010",
      "010001101001101000111011100101",
      "110011110100001001110000100000",
      "010010101001001110010111100001",
      "110111001101111000011101101110",
      "000110010110111111111001010111",
      "100011000111010011110001100000",
      "000010110101011110110101010101",
      "001110000110101110001100010001",
      "000010000111100011111110010011",
      "101011011000110110101001000110",
      "110011011001110001100001001111",
      "011110100101000010010011000000",
      "110111010011101100001110100111",
      "010100001110001110110000000000",
      "101110110001000011111011101001",
      "100111100111100001000010000110",
      "101001101101100101001111000011",
      "100001000111001110011101011101",
      "110101110000101110011011100001",
      "000010011001101010101111011000",
      "111100010000101000111000110100",
      "000100110101001110011110010001",
      "000001000001010011010100000110",
      "011010011010100000000111011100",
      "000111100101100111000110110001",
      "111011101100110011110001001101",
      "101101100010011000011011101101",
      "011011101011111010100000011001",
      "001001100000110110110100111101",
      "101010011001010101110000011000"
    ),
    (
      "011010101111100100101010000000",
      "101011000101011111110110110100",
      "000101000111010000000110011111",
      "010000001011110110111000010000",
      "110011111100111111111110010011",
      "100010011000111111000100101000",
      "010101110111010010111000000001",
      "111001111001011111110011001110",
      "111101001010111111110001010001",
      "100010001101110111100100111111",
      "010001010010110001000000101001",
      "010011110000101010000100101011",
      "011000111101001011100101101100",
      "101010001000011111011010101000",
      "110001001111101111010111010111",
      "110011111000110111110111010111",
      "111111111001001000100000110001",
      "101011111101000110011110111100",
      "011001001010101001001010000100",
      "001111001100110010001111110101",
      "011000001100000100011010011100",
      "010111000101100111000110111010",
      "010010100111010011000110111111",
      "001100110110101110100111101100",
      "111101010101101000101101011100",
      "011110111101111111101001011000",
      "011111010001000000100100011000",
      "100110100110001110010011111101",
      "111000001101011010000000001011",
      "110111011110100110100100000110",
      "110111000001011111111100011010",
      "010100001010000001100111101001",
      "001111010011000110010011011010",
      "101001000101000110001101000011",
      "111110110011000001000001011101",
      "010001101110010110111111001000",
      "011011010001011010101010010000",
      "001110010100010011100111000111",
      "100001010100011001000101110001",
      "110110101101011110001000001001",
      "110000000111110111101100001111",
      "101000100110111100101001101000",
      "111011001010011110110010011110",
      "100111110110000100111111101101",
      "101101000000000100100110010110",
      "011110001110100010101100000100",
      "111110010111110101111111000101",
      "111100010111110111010010001001",
      "010110001011000100000101001110",
      "100001111011010010110111010010",
      "001111100100001100100111110010",
      "111110001111100110101110101111",
      "100110101111010111100000101101",
      "100100000111010010011010111101",
      "001100011001110101001011010001",
      "001100000011110000100001001101",
      "101011101100111100111000110001",
      "111000011111111000000011010110",
      "110110100010101100110011100010",
      "111110110001001111001001010101",
      "001101111001110111010111101111",
      "111110011001011111111010001110",
      "111100100110100101110010000101",
      "100011101110110010000101001110",
      "111011000010100010010010111011",
      "101111101110010010101110101011",
      "101011011011101100010000000100",
      "011110001100110001101110110101",
      "100010000000101001000100010000",
      "110011011010101011011001101001",
      "100100100110100000011011100001",
      "111011010011010101100000001101",
      "111010111010100011110000111000",
      "100101000111100101001000010010",
      "110100011111000001001011111100",
      "010110110110001010100100011100",
      "010001010100101010010010101010",
      "101001000101000110000011100010",
      "111100101000000101100011100111",
      "101111100001101101100001000111",
      "110010110101000010101100111011",
      "011011111011000101000100011110",
      "110001101100100010001110010000",
      "100010101000100011110101111111",
      "010110010010111101101111010101",
      "010101011110010111111010010011",
      "100101101000100101111101110000",
      "100001110110000100111000011111",
      "101011100001010110100111100001",
      "101000010011110000011001001001",
      "011110110100110011001011000000",
      "001110000110100000011100110001",
      "010001001001010110001000111100",
      "110100011010001010000110100100",
      "011011010010100111110100001010",
      "100010010100101000101001011010",
      "110011111000110010101111101100",
      "000010111110001101111110100100"
    ),
    (
      "000010011111101101000011101100",
      "111111010010110000110101001011",
      "100111110101110000011111100010",
      "100000111110010000001011001101",
      "000101100011000010111101011110",
      "000001011000000000001000101100",
      "001100111010101101111100101111",
      "000101001110100101101110000010",
      "000001100010000000000100010110",
      "110110111100110111001001000000",
      "011000101001101101000010010011",
      "100000111011000100110000111110",
      "111101001010111010110011101001",
      "000101100001010101110100011110",
      "111100111011100010000101001101",
      "001010110110001010110011010011",
      "110101011001111010101010011111",
      "110111110101000101001011011000",
      "101001100100111000000000000111",
      "101010100010010100110100101100",
      "101010110100011110100110000010",
      "000111111001011100001000110010",
      "001001001000011101000000000000",
      "110101010111010001001001000100",
      "000110111011001100010011011100",
      "010100100000011100011010111000",
      "010011110001101011110101011101",
      "110110110001110001110011111000",
      "010000111011110100111010000010",
      "101100101010001110011101010111",
      "111111000000110001110110101011",
      "101111010001100100011101001100",
      "001010010011110111001101100111",
      "110011111110110000101100010110",
      "100111011001110001100000101010",
      "101011111011110011011000101000",
      "000100001001110111001110010100",
      "111110100011100001011000111011",
      "000110100001101011110111111111",
      "100010110110010101101100001010",
      "000110101110000100001001111001",
      "100100101101000111001000010111",
      "010001001010000101101001001110",
      "001100001100101111001100111000",
      "011100111111111011101101111110",
      "001000000001110100011101011111",
      "010111011001110000110011001001",
      "010111111010001101110111011010",
      "111100110000110001100010110101",
      "100001001010000100111101000110",
      "010111011010111000000101100100",
      "011000110011010110100110011000",
      "001110110001111001001000011101",
      "110100001101011111110001111001",
      "000110101000101001100101111111",
      "011101001101111111101010111000",
      "010010001011010110010001110011",
      "111000110001100101110110000110",
      "000110100011001111001110101000",
      "001010111011101111001000110011",
      "000111001110100001001011111110",
      "111110110100110100110101000111",
      "001100111101010101101101011100",
      "001100011001100110101110101111",
      "000111111011100000011010101101",
      "101100111101100000101000011001",
      "000011010111001011111011011011",
      "100001101111110001101011110010",
      "111000011011101000100110111001",
      "100110010001011111101110111001",
      "111111011011100100011110001010",
      "110111100110111100111011111110",
      "110000100101100000010011010100",
      "010011001110001001111011000000",
      "111100011011110110100010110001",
      "101000101101001011001010101101",
      "001001010110011100101010001111",
      "000011000010001100100010111101",
      "100001011010000100111000110101",
      "110111001010010110100110011100",
      "011011110011000000101100010010",
      "010010010101100110101010011011",
      "010100110000101010100011111101",
      "111010111101101101100101101110",
      "101011001101001101101101110100",
      "101111011100111111110000000000",
      "010001010010000010001001101100",
      "001011100100101110000111001010",
      "100101100100100100010111010000",
      "111111111100010001100110101110",
      "000101010100011110100010111111",
      "101101001110101011000010001101",
      "100111111000101011110101111011",
      "111100011011000101010011111101",
      "101110001101101000110101101000",
      "100000101000000000100111011111",
      "110011110010110101101000011111",
      "110101100011101100111101001111"
    ),
    (
      "000100110000111101111110001011",
      "001101110000011011100000100111",
      "001110010011001111000000001101",
      "100111110101010011010110100010",
      "000010011000001111010000000111",
      "011000001000011010011011001111",
      "100100001100111011110101010010",
      "000101001111011111101101001001",
      "100000101100001001101111011000",
      "001001101101000100100110110100",
      "001001101010100100001000111001",
      "111110101010011100110100101100",
      "001100111000001111000010111101",
      "111000110001111000110000011111",
      "011111000011111001110011100010",
      "100000000011011100101000000101",
      "111010111011011111100010110000",
      "000010000010000101100111101110",
      "001111111100101010000011111011",
      "110110110000010011101100000101",
      "101001111001101110000001110110",
      "101101010001001010001100010001",
      "111011111001111001011011100000",
      "000010111000011100001001011111",
      "110100100100001101110001101001",
      "001000001011000010001001111101",
      "111101001101100101100011000110",
      "100001001101000001010010100010",
      "110000100101001111101001000101",
      "101001111010101100010011001000",
      "100001000011111111101011101110",
      "100111100111000001100101010010",
      "000010111001110100010101101110",
      "111000110100100001010010111101",
      "110011011000010010011101000011",
      "100001111011001000100100001110",
      "001111010100010111101111101111",
      "111101001000001110100011100010",
      "010010101011110101000101100010",
      "101000011111000101100001010111",
      "000000010001111010101001110010",
      "000000101011111001001001010001",
      "101010010111011111000101011001",
      "110110001110110000100000110111",
      "101010110011011011001100011101",
      "100111101001111101110000001101",
      "000100100101100011101100011001",
      "000111010001111011010101010110",
      "000111111101011100101001000011",
      "000100011001001110111000101101",
      "001110101111011110111000011100",
      "101000110000101010001000010011",
      "010111001010111100000001110000",
      "110000101110010100000000101100",
      "000101010001110001011010000010",
      "101101001110010011110110110111",
      "111101010110010101010011111111",
      "100101110100110001000100010001",
      "000111000101111100001011001110",
      "011000001011010111001011111110",
      "111101001001100011101111010110",
      "110101010110000011100011000101",
      "001101100011111100010101011110",
      "111110001000001110110000111111",
      "001001101011101010110110001110",
      "001000101011110011001100101110",
      "000010111010001110101101101101",
      "010110101100011110000001100101",
      "001010111101000010001111110000",
      "010001110101111000010010100001",
      "101010111011011101111100000000",
      "101010111110000010010000100111",
      "011001001100100010110010011001",
      "100101011110000001000001111011",
      "011001111110101011111010101111",
      "110000111000001110100111000011",
      "001000110111001111100010000101",
      "100000100110110101110010011010",
      "011011111110000100101111000011",
      "111010011101011111101110101110",
      "100101110110010110000010101000",
      "111100111000101010111011111100",
      "100011000111010110101111001010",
      "111011001101101011100011000011",
      "110111010000010011000001100101",
      "011111111001101001011010101100",
      "001010010010010111111011011011",
      "001010111001111110100101000110",
      "011000010101101100011011111110",
      "110110001010011101001111101001",
      "101010100111000010010010011110",
      "011101111010101000111011000011",
      "010001000100101110010010000111",
      "101110000100001110101101011110",
      "011111001010001000100010001100",
      "011111111000110010100111001110",
      "101101110100000100000111000100",
      "000101111011110011111100010000"
    ),
    (
      "111110101011110001110011101100",
      "000100100110110000100110010110",
      "100101111110100010101000110101",
      "100000000100010001110111011001",
      "010001100110110010000010111011",
      "110000101010010001110001110100",
      "100110100111111110000100011100",
      "110100100100000110111010000111",
      "110001111100101101000101110011",
      "001111111100001000010110101100",
      "001010111010000101011111000010",
      "101101000010011111100100110100",
      "000101100010111111100101111101",
      "110010010110100001100010110001",
      "011110000010011011001000011010",
      "110101000111110011011010101100",
      "001101011110001110000011111011",
      "001111010000000011110011100110",
      "101001010100001111010110110111",
      "110010111110011100111101100000",
      "011100111111010011111100110100",
      "111001110010101100100001001111",
      "111110101011110111101010110001",
      "011111011111110001000000011100",
      "000110100000111101001101110101",
      "100101100001001010010101000001",
      "010111000011111110001111111100",
      "010010001001111101001011000100",
      "000110101011100101110110101011",
      "110101000000111111101101011010",
      "001011101101001101000111000001",
      "001000110110000010111100010101",
      "100111011110001001000111100101",
      "111010110000001010100010010101",
      "010010110111011000010000111100",
      "111110000100111100011101011000",
      "111000111100100011001101011000",
      "101111010010110010100000000110",
      "111010110010001011100011101011",
      "000111001110011101100101111111",
      "110100111111101001100001000111",
      "111101000111111110001011111111",
      "001010011111000111001000011011",
      "100000110001100011110101001001",
      "011101000110100001100100010010",
      "010100101000000101100010100100",
      "011100100010100000110001001011",
      "011111001011111111011101101001",
      "101011001100010010100001000101",
      "001100001111000000000001101101",
      "100010110110011010111011100110",
      "110011101111100101000110110001",
      "100101111100001110101101100111",
      "010100111001010101000001100000",
      "100111110000100011001000010110",
      "110111110001011100001101101001",
      "100001000111110111011110010010",
      "011110010010010110110001101011",
      "001001101100010000100001101100",
      "111001101010101010000110010011",
      "011011111000010000111101100111",
      "010001100111010101001000100100",
      "101101100101100110000011001011",
      "110011100100101101100111000001",
      "111101001000001111010110101101",
      "111010111100100001111110101001",
      "001000101011110100001011110111",
      "111111011101110001110100001000",
      "111000101001000001100111001001",
      "000010001001111110000010001100",
      "100010010000001100000111010100",
      "111010010011000011111001111111",
      "101100100100011001101101000110",
      "111111011101100101111110110000",
      "000011011110100011010010000111",
      "100110001111111010111000000111",
      "111101110000010110101111110001",
      "010010110110001001011111010110",
      "111010100111110000010011100110",
      "100010101000010111111111001110",
      "001111000100100101011011010001",
      "011111101110101001000110100110",
      "010011100101100101000011011000",
      "111000100011011111000000011100",
      "110100010001101100010010011110",
      "110101001010010010011100000111",
      "101011110010010011001001110100",
      "110111100110100100101111000111",
      "010010111101000101001001111001",
      "110100000110110111000001110000",
      "000101100001010100101011000100",
      "000101110101000000011001100010",
      "000100100110101110100110011011",
      "000101111011111010100111111011",
      "001000111011100010010100100100",
      "001011000000100100001000101100",
      "011100000111101010010011011000",
      "000000101001011111111100011101"
    ),
    (
      "011101011101000001101011001100",
      "010011111010011100111110010000",
      "010010100011000110011111011010",
      "100111001111101010110011001101",
      "011001000011100111110110101100",
      "100101101100011010001001111100",
      "110111101010010100111010011111",
      "000001101001000010110000001011",
      "110011101110001001010000010011",
      "001001011101110010000111110100",
      "010010110011000001011100011111",
      "100100000011000011011010110110",
      "011100010111111111111111000000",
      "001011100000001100001000110101",
      "011111000001000100111101110110",
      "100101011011111000000001100100",
      "100100000011110111100101000100",
      "011010101000011110111010111010",
      "110011101110011101000110010110",
      "111010000010111011111001011001",
      "110111100001110011111010001110",
      "011000100001000011000110000011",
      "111010011111010101101111111000",
      "011000101100101100011011010101",
      "110000110010000110010000111010",
      "101000001000000000011010011101",
      "110110100111101010110101101111",
      "110111001101110010001111110010",
      "000001111110001100011000101100",
      "101110110111001110010100011101",
      "000110101111000000111111100100",
      "100100000111001001110101010001",
      "101100011101011000110100011000",
      "101011101011111101000000100100",
      "010100010111101010101101010100",
      "111111110111000101000110011110",
      "101100011010110100100010011100",
      "000000100001110100011101011111",
      "000110010010001110000000110101",
      "001110011010011010011111100101",
      "101001111001100000100101001101",
      "011101110110111110100100000010",
      "101001011100011010101111111000",
      "010001011000010010010011011100",
      "111011100010110110111001000000",
      "111101100111100100110111111010",
      "011100001000000110110010000001",
      "111001010111000110110001110101",
      "101111100001110011100111010011",
      "111101000010001010001111011110",
      "010001101110110001010001011010",
      "101010001100000011001000100000",
      "111011001110000111010001110111",
      "011101101010000010101111011100",
      "110011111111001001101010100011",
      "000010100111101100011000000010",
      "111000010000100001010010100110",
      "010001000001010011110001010011",
      "010000001001001111011000001101",
      "011001111001001011011000100010",
      "110001010011011110001010010100",
      "010010001110110101001001001010",
      "111011110001110100010100001011",
      "111011011101010001100110000100",
      "100001100001000010010100001100",
      "110101101111001011111101110011",
      "010110101100011010011111111100",
      "111001001001011110100100000111",
      "001111001000001110010101000110",
      "100111100111000101010100010101",
      "111001010001100010010011101000",
      "101010111110010010001001010100",
      "110011100110010011000110100010",
      "000111010101001001011100111011",
      "101000000001111111010001011110",
      "010110101100101000011010101001",
      "101011000101111100111110011101",
      "001010100100110011100111111101",
      "000101011110010001001001101110",
      "010010010000000101000000110011",
      "111110111010100110100000001111",
      "101110111110111010101011010110",
      "000011110111011000110000110011",
      "101100100000110001101100011010",
      "111110010101010101111001110010",
      "101110100100000010111010010101",
      "101110100001001110011111000111",
      "001101100000010001010111111010",
      "001111101111010000101000111110",
      "110011111001011111110011110010",
      "010000110111111100001100111011",
      "100111110011000011000101010011",
      "000011001000111100101101010101",
      "000101100110110110001000011111",
      "000000010110100001110111110001",
      "010000011111101101010101101110",
      "000011000010100100111001000001",
      "101010110001010001011000011110"
    ),
    (
      "111011111011010011110010011100",
      "100001100001100001101001011101",
      "001110001110110000000110010101",
      "010000011110110110110000001001",
      "111001111001001111101100001100",
      "011001000100000110010001101100",
      "111000010110100100101011011111",
      "001101100100110110010111001101",
      "100001001010101100110110110101",
      "010111001100101110100011010001",
      "110101111011000111010011111000",
      "001010010011001111101000010110",
      "110001111100110100101011000111",
      "011100110010100111001001010110",
      "101100010111001000100000111110",
      "000100001101100110011111011100",
      "011101011100100101011011101111",
      "100100001111011000110010000101",
      "000110010100001110001110000111",
      "110010000111111101011111100001",
      "110000100110011010011101101111",
      "010000101000000011000100010001",
      "100010111001000001101110011011",
      "111001100001000100111110101111",
      "101011010110011000101111010111",
      "011001111001101111010001001111",
      "000110100000010010101110101010",
      "111001111101101011101011011011",
      "000010011001010001000001110110",
      "110001010010100010101011100011",
      "000101001101000101100101001011",
      "011100111101110100001111010010",
      "001101110100001001110000000011",
      "101000110000100101010001011001",
      "001110011111010111110011110001",
      "110101101101010001101001101101",
      "100010111010000111000000001111",
      "010000000000111000100100101011",
      "100111011001000011100000101111",
      "111111011010010011011101110011",
      "010101110100100101111101111001",
      "010000001010111100011010000011",
      "000111011110100110100010010100",
      "001101101010100100000110101101",
      "100000100101100010101111010010",
      "100100000100100011100001010010",
      "010010000001110000111011011111",
      "100010000110001000010001000111",
      "101100110110101111110101111011",
      "110010001101010110001111010100",
      "110010101101010111000001010010",
      "000010000000011110000101010100",
      "010011000111001000110001010100",
      "001000111011011110001000111111",
      "111110001011001001111111101110",
      "111000110011111000000100110101",
      "010001110011010100101010001101",
      "011100101111100101101001010011",
      "011001000000111101000101111101",
      "100101011010100001011110011111",
      "011111110001000001111000011110",
      "101110101010010111000011110111",
      "001011011011001110101000010101",
      "000001010011011011100010011010",
      "111010010101010111101000010100",
      "000101101001100011000101110000",
      "011010100000100101011100001011",
      "111010001011100111011010011111",
      "011011101100110001010110110011",
      "001001011111101111100111111000",
      "010110101010000010111101110000",
      "001000000000010010010000111011",
      "011110101011010011010001011000",
      "010000100010010001001111111001",
      "111110110101000111101110100001",
      "011001010100001101100110011101",
      "100111100000111010111101100010",
      "011100011011100011000111100110",
      "100001111010001110101010110110",
      "010111111100110001111001001011",
      "001100000100100101010110000011",
      "011110000111011100001011100110",
      "111111101111000111110001010101",
      "000110001010100101111010011100",
      "001110101011011000011111000111",
      "101111001100100011000111011111",
      "110110010101110101011110001110",
      "000011111101110111000001110010",
      "000010001101111110111011011010",
      "010101000011010100000100111011",
      "011100010010000000001001001000",
      "011000110011101101010010010111",
      "100000001100100100110101110001",
      "110111011011010000110110011001",
      "111011101011010000111110100110",
      "000101011001111000000001101010",
      "110000010110010110011100110100",
      "010101001100100100110101010011"
    ),
    (
      "010000101100000101100111100010",
      "100111110001000010111010001110",
      "111000111111111111010110001101",
      "110111010110101100010011110100",
      "101101101111111101001110001100",
      "010111111011000010011110011111",
      "010001011001011001011001010010",
      "000110001011110100100010110010",
      "001111111001100001011000000101",
      "000001111110000010110101001011",
      "000111001000011101000110000100",
      "011111111100100110011101000011",
      "111000111101001111111101111001",
      "111110000111101111011111001000",
      "101000000011010011111100111110",
      "000010001011111111000000001100",
      "101011101100000000110011100001",
      "000110100100101000110001111001",
      "100111010101101101111010001010",
      "010110100111001011100001011001",
      "111011110000011111111001000100",
      "001101100110010100101100011010",
      "110011100011011100000011111011",
      "101001011110101101100101011101",
      "001110110011000000110001010101",
      "010101100101100011010011011101",
      "010101011001111110111001110011",
      "010111101101010011101100100111",
      "010001110001101110000000110001",
      "000100101010101101101111001000",
      "111100010011000111000100010001",
      "000110010100101011000000010011",
      "010110000000010011001011011000",
      "110001011111010111000000011100",
      "001101000010100000000100001111",
      "011000100111110100010110011000",
      "101010100001110010000010000010",
      "110010001001010001100000100010",
      "110000001111000111001001000001",
      "001110010100011111001111011001",
      "101110000001001101011100000100",
      "000101000111000101100110010111",
      "101001010001011010000001001100",
      "111000000111011100000101110101",
      "110100001000110110100001010101",
      "001001100011001100101010000011",
      "011100011010100101011011001010",
      "100011110001101001110000101010",
      "001010001010010000010001010011",
      "010010001010001001000011001000",
      "111010100101101011000001000010",
      "111001010011110000011111101111",
      "011101100011100001110101100010",
      "000110000111111111101010011100",
      "000010001001100101111001010000",
      "010101101110010011101110110000",
      "101100100111010101001110000010",
      "110111010000110111101110111101",
      "011100000010100000111000011001",
      "111010100111100100011010111110",
      "111001111111011010111110101010",
      "011001000000000001000000000110",
      "100101001001011011100101011101",
      "011100011101101101100011111101",
      "010110010011001101111101011110",
      "001110110111010110100001000010",
      "100100111010000100101010111100",
      "000011011000100011001100101100",
      "111011101100011101011100011011",
      "011010000110110111111111001001",
      "011010001011000101000100101100",
      "111110001000001010001101110100",
      "100001110100111011011010000111",
      "101110001111010001110101101001",
      "011010100000110110100010011100",
      "011110010111100101101111100110",
      "011111100101100100111001011110",
      "001011010011111000110011010101",
      "110000111011010100100001100010",
      "001000001100000111100011101111",
      "110111010000101111011011010011",
      "000100110111010001011001011001",
      "111100110010000110111011101100",
      "111001101011111110110010011100",
      "000001011110011000001110010011",
      "110111100001100011010000011111",
      "101001111101101101000010011011",
      "011111111001111001100111101100",
      "110001010011101110000001011110",
      "001000011100111110011111110001",
      "011011110010101011111100011100",
      "011100011111000111001101011000",
      "001010101001111110110010011010",
      "100000111111001111001101000000",
      "111100011111101011000000101110",
      "010100111101011111000011000000",
      "000100101011100011010011000100",
      "100011111111111111101100111010"
    ),
    (
      "001110101110000001100001111000",
      "001101100000000101110100011100",
      "101110111010011010010000101010",
      "110010111100101010011101000001",
      "101100110100010101111100000010",
      "110000010000101111101011000011",
      "101100011000100100010001101001",
      "001100110000001110010000111100",
      "111011011101100101010100100000",
      "011010010101000101000111100001",
      "111011011011011101101001110110",
      "111100100000010100110111011001",
      "101000101010000110101100001101",
      "011101001100100101011011100011",
      "110101000110010011100100001000",
      "001101000110001010011111101001",
      "111110011111101000010100101010",
      "110000110101101111100100011001",
      "010101011000001101010010100111",
      "000011100110101100010011000111",
      "001110001011010011100100011001",
      "000110110010101101000100000011",
      "011111011100100110010100010110",
      "101001001001001111110110011110",
      "010001010010101111001110010001",
      "101111000111110001010010000100",
      "110000011111100011100111100111",
      "011001000100000000110000110000",
      "001111100010001001100100111111",
      "001111000010010000111110001001",
      "000010111010110100111000011000",
      "010010000110011011011111101100",
      "100000111110010111110010111011",
      "100000100001101100001011000101",
      "110010111010001111010010100111",
      "110001011100000110001001111101",
      "001101100000100111101100100001",
      "111001000100110100101100110100",
      "011010001111000100111011010011",
      "101000100000110000010001111101",
      "110001101001100011111111111011",
      "111100111101100101011010001111",
      "001101111110001111110111000001",
      "010001100111110101111010011101",
      "000010010111111101001010111001",
      "110100001011100001101111010100",
      "111010110111110100100100100110",
      "101000111010100111100110001000",
      "110001010110011110000001110101",
      "010000101010110010000100000010",
      "000100000100000011001110111000",
      "010000100001110000001111001001",
      "011010001011101010010101110111",
      "011011001101010110100011010101",
      "010010000110101010100011110011",
      "010110100001101100010010110011",
      "111100111101101000010101110011",
      "010010011000011000111111110101",
      "011100110111000110001010100101",
      "010000100001101111100000101100",
      "010110111001100101110000011001",
      "010011001110101011000110100001",
      "100011011001001110101100100000",
      "011111001000111011000101001011",
      "111111001101000111100000111100",
      "110011011100001110101000011110",
      "110110111110001000001001101110",
      "010101001101011100111001001110",
      "110000100011100110001010011010",
      "010101101111110101111001001011",
      "110001101000101000010011000000",
      "110010101101001100011111000101",
      "110011110011101000100011111011",
      "001011101101001101011010000011",
      "011111111100010011011111110110",
      "011001010110000101010100111001",
      "100110111100110110101001011101",
      "011000010011010100011010111100",
      "011011001111000111011010110111",
      "100010110011101000101010011100",
      "010001111101110010001010010110",
      "011101101001000001000010101000",
      "100000111110111010110001110101",
      "100000001011101100011000000010",
      "000011001000100101010001100000",
      "111100111000110101100011010011",
      "111110110100100101101000110100",
      "110111000001011111011001010011",
      "000010010001101001011001010011",
      "000111011011110011110011011010",
      "110000001111101110110001000011",
      "101010100011111110010011111111",
      "101110011011011010101111110101",
      "111100001001011111101001111101",
      "011101010111110100101011100010",
      "110010001011100100101010010100",
      "110010100111110110010100010101",
      "111001111101001001001010110000"
    ),
    (
      "001001111000110111011000011110",
      "001101101100101101010101101101",
      "101110100100111000110000100011",
      "111100001001011101101001000110",
      "010101101110110111110011000000",
      "101110111100100111001001100100",
      "101001110100101011111101010011",
      "101000000111101010010011101111",
      "011010001000111010101010110000",
      "000111010100000011100101111111",
      "111100100011011111110110010010",
      "110110110011111100110100010111",
      "011010001110110011100010101111",
      "110110001000111110110100100011",
      "110011101011110000001000001000",
      "111000100010011001010011011100",
      "111010111101101111111100000100",
      "101110000100101000000111111010",
      "001001100110001010100011001001",
      "010010000100000011101010100010",
      "110010101110110100001110011100",
      "101110001011000010111000101001",
      "001100000011001111000101010111",
      "011001110100001100100100000110",
      "101001011110011000100011101001",
      "010100011011001010000001000000",
      "000001010101100000010011000101",
      "100010101110001100110100111001",
      "111101110001100000011111111010",
      "011011111111110101100100110110",
      "001011110100000000111000100011",
      "000100110100011101111111101100",
      "001111100011010010011101001011",
      "011001000010000001001100101101",
      "110100101010000100111100010010",
      "101000111000000100110001010011",
      "001110010110110111011110111011",
      "110001111111111000000010100110",
      "111101011011101100110011011010",
      "101010001110000001011001101100",
      "101101110010011010110110100010",
      "110110011110001111000111000001",
      "010001111000110100110011001010",
      "100011001000111111011101100111",
      "111000011000010000000101101111",
      "111011100101010011010011000100",
      "100010001100011010010100000001",
      "111101011101111001011010111001",
      "111101011111101010000011010010",
      "111011111011111010111110101101",
      "101111111010000110001110011111",
      "011100101010010010000010101011",
      "100100110110110111100011100101",
      "001100000010100000111001100010",
      "000000011011110001010001010000",
      "011001110000011010010010111001",
      "100001001111110111101011000001",
      "101010111010001100000011011011",
      "011100101101010011001111000101",
      "110111011010101111100111011101",
      "011000010011010101101001110010",
      "111001110000111110100011101010",
      "100011110000010100001011100000",
      "000000101111010100011111001111",
      "011100110101110110010101110110",
      "011011011010110101111100010011",
      "011010010101100001000110001010",
      "110100101000101101001011000100",
      "110010101010111100110000001011",
      "011110010111101000110111010111",
      "110101111001100110000010000110",
      "010100011001001110101101010010",
      "000100100110011011001000111100",
      "100011100011000010010000111000",
      "001000011010000001010100011010",
      "011100101001111110111010110100",
      "100101110000110010111001111111",
      "011000000100001100110110011011",
      "010100011101101001010111010001",
      "110010100001011111000110111011",
      "110100010011011001000011100101",
      "001101101000101101011110110010",
      "011100101100100101100111011010",
      "011010000001000001111010110000",
      "101100011110110110010011100011",
      "010000000101110001000001111111",
      "000010000010110110010001100110",
      "101011101110100100110010010000",
      "100010100010110111000100110101",
      "100010011111110011010111111101",
      "100111011110001111010000010001",
      "100011011010110101111111100110",
      "101000100001001011001111010001",
      "100010110010100000011010111100",
      "010110111111101110111001111100",
      "101001011100101001001110100101",
      "011000101111010110101011001000",
      "111101001110100111000001011000"
    ),
    (
      "000111010000001000000010100000",
      "000000011101001111001001100011",
      "011010001111111011010100010001",
      "010010000000110000100011001100",
      "110000110001011010110111011101",
      "101010110100010111111000110100",
      "001001111111100111011010111001",
      "111011011001111100111000011100",
      "110110101010010000101011111000",
      "110101010101101111010011110110",
      "011101001100100000101111001000",
      "101100101101101110101010010011",
      "101001011101000010010000100111",
      "000000101100110010011110010101",
      "011010010000011000010001101011",
      "101110101010010000101100111011",
      "101110000010001001111110101111",
      "011111110011110001111011000011",
      "101011100011001100110110000000",
      "111011000001010100001011101100",
      "011011101001101001001001011111",
      "101000110111110001111001000011",
      "010010101000110010110000101001",
      "110001001010111110101001011110",
      "010110111000111010010111010000",
      "101010101101011010001110101110",
      "100100101011010000001100000000",
      "101001010111100110110000101011",
      "010011010010110111001110101101",
      "100101000100110100110010000010",
      "001001000000010001001000001010",
      "011001110011000100010010110101",
      "101110101010111000100101000001",
      "111001000010001010110000101000",
      "000011011011001010111111010110",
      "100000011100001101100000101011",
      "101000000101110011101110110000",
      "101111101100010000000010001100",
      "101000110001001010101011010010",
      "110000100110000011010100011100",
      "000100001011001011101010111001",
      "001100111001000111101000100010",
      "001001101101100010001001011001",
      "101100101011010100000011001000",
      "001010000001100001001110010000",
      "111110101000000000000111101111",
      "011000001001100011101000100010",
      "101000000100100100000110010011",
      "101101010111010000110001110000",
      "110110000011100000001111010101",
      "001111110001001100101001110001",
      "010111111110011111011100110010",
      "011010101111110010000001000110",
      "101110100010101111100010011001",
      "010000010111011000111000000001",
      "001010001101100011110011011000",
      "110000110111010101111000001011",
      "101000000011100111110110001011",
      "001110110000110110111011000000",
      "001011100111001000010001011111",
      "000110010101000010101101101101",
      "101010000110010011100100000010",
      "110001010001100111111101100010",
      "100000001000110010001100110010",
      "011111110010000001001011000010",
      "001010101101010111100011001101",
      "111011100111100100110011011010",
      "110100001001100101000110011000",
      "010111100011111100100000010001",
      "100110010000011001101101100111",
      "010110100001100001100010110001",
      "001001101001101000001001101110",
      "110101000100111011011110111010",
      "000111011001011100100100000111",
      "100110100011111111100000011001",
      "010100110000110100000001000110",
      "110011011110110100011100011111",
      "010111011010100111000111100010",
      "100110110001010100101101011011",
      "000011011010001001110111110101",
      "111101011101010000101100101100",
      "111101011111110110011100000101",
      "101010110001001101000111011110",
      "100010000110100000011011011111",
      "001110000100100001001100000100",
      "101110111100111101101001111000",
      "101100001000011110010110010111",
      "110100011010100010010001100001",
      "000100011101001010011010001101",
      "111011001001111001010110000101",
      "011000000100101111000001000011",
      "100010110110010011110011111001",
      "011011101100010001111011110000",
      "011110010111101100101111110011",
      "111110010000000111100000000011",
      "111000111001110100000110100011",
      "100011010001110100101101000000",
      "000100110011110001011001100010"
    ),
    (
      "111001000011000010001101111010",
      "000111000000110100011000011010",
      "011011010111010101010101110001",
      "101111010101000010100001000101",
      "110110111010110001100111100111",
      "001011100001111100000111100011",
      "000111100100111110000000100111",
      "001100000010011101011011111111",
      "010011000100011101111111000011",
      "110000000100111000111111111100",
      "111101100101101011000011000001",
      "011001100001101100000111110010",
      "101101101111010111011110101010",
      "010111110011011010010001000010",
      "010010010001010001011010101100",
      "101000001011110011100001100101",
      "101000011111101010001111001010",
      "011111111101010011111111010111",
      "000001110110011111010011101000",
      "101111011000101100110100111010",
      "100010100010101101001011110011",
      "100111100101111100101100110101",
      "000101001001010011100011000001",
      "001101111111111000010010011010",
      "010010110010011101100001010000",
      "101111010101110100010011001111",
      "000111001001100001010101010011",
      "000001100001001111110010100100",
      "110000111110111000100100110011",
      "010100000000101100110001110001",
      "101101111000111111000110011110",
      "110101100010100000100001111111",
      "111101010100011111011100101010",
      "100111001001101111001100000101",
      "111011000100010010101010011111",
      "101001111101011111101010000110",
      "000100101000000111000011110010",
      "101000111000010111110011000010",
      "000101100110110010101010110111",
      "000101001000100001110000110100",
      "100100010000101010011110111010",
      "100000011000110000000011000101",
      "010111111100100110111000111001",
      "100011101100001110000000111011",
      "011001101100101011101101001011",
      "111000110010111010111000100011",
      "010101110001110101001011011011",
      "111010100100000001001101001101",
      "100011100010001011111111010101",
      "001110101000101100100101111110",
      "111101100011100011000101110001",
      "011010000001111001011011000100",
      "010011100110001010000110011101",
      "110010010001100100111010101001",
      "001101011000100011100011000111",
      "000110101001010001111000000110",
      "101010110111010110100110101101",
      "100101101110000101111000110000",
      "000000100101111010001110000110",
      "001101101011000010101101010001",
      "101101010011000001010110001110",
      "001011101001001100101010110011",
      "101011001111011110100010110100",
      "101111111001001110100101101111",
      "001010001101010101010000010001",
      "100110010110111010101011110010",
      "111110010011110001000100000010",
      "100011010101101110010010010001",
      "011110000001111100100110100011",
      "011111111110011010101111110010",
      "101110001011111110110100100011",
      "110101110101001010000101011101",
      "100001011000110000100001101100",
      "110111110000011111011000011011",
      "001100001110001010001100001010",
      "111001111001100000011110000101",
      "100010011101000010011000101010",
      "000011100100000001001000001001",
      "011101110110010100001001101000",
      "111011010000101110011100001001",
      "010011111000000000010000000110",
      "011011100100101100001000001111",
      "000101011111101011100110111000",
      "000010100111001001100001010010",
      "011011110100001110101001110011",
      "100110010001011111001000111101",
      "011001000101100101100100001111",
      "011000011011001101000110110111",
      "010010011101001001110001000110",
      "001001000011011001100011110010",
      "100100001010010110000101111111",
      "100111111001010111001101111010",
      "100111101111101101010010001101",
      "011110110101011000011110101011",
      "010011100111000000011100000011",
      "101001110010100111111001010001",
      "100101001111110100100111101110",
      "000100000001110101000100001101"
    ),
    (
      "001110111100000000011011100111",
      "111101111001011100100011010010",
      "000001001111110010111111001110",
      "101110000000101101010001011101",
      "111111111001010010000011100010",
      "011100110001110111110100010010",
      "000001011011101101110100011100",
      "101100010101011011100100000010",
      "001000110100100011001011001011",
      "110100010100101011001000010001",
      "100001001100000010010101011101",
      "011000010111010010010000110000",
      "111101110000000101001000000001",
      "110100011000011111001101011001",
      "110010110111101101010011110011",
      "010010110010111111110101110011",
      "110001000001111111101110101110",
      "010100010000111000001111111001",
      "010011010111110110010000010101",
      "001000110000010011101110001010",
      "000100000011101001011100111110",
      "010000000010010000011010101001",
      "101001000000101010101011100100",
      "010010011111100011001001110110",
      "011011101111011111011110101111",
      "010010001000110001100100011110",
      "000111101000100111011010001110",
      "101001011101011011100111011011",
      "010100000100011111110110010010",
      "111100101000110100001100010011",
      "101101100111100010011000101110",
      "100000110110000001100000000101",
      "010010110011110111100010001111",
      "000010001101100100111100110001",
      "100101010100011001000011000001",
      "101100111000100110111101010101",
      "000110111101001101110000011100",
      "110111101000000010100110110011",
      "100100110010001100100101111100",
      "011101110101001111011101111110",
      "110000000010010101000110101100",
      "100010110001111011101000101001",
      "110010011101011000110011010101",
      "100010001011010010110000010101",
      "110100110010011100101100000001",
      "000110110010100110011000001001",
      "101100001000001010100000111001",
      "011110001110100110001010111010",
      "111000111110001111110110101110",
      "001111011111000001000001010111",
      "101011110001111100100001111100",
      "101000001001100010101010000100",
      "010011110100111000100000011110",
      "100010101011100001100101101000",
      "111101010100111001100111101111",
      "111011000010111001110110011100",
      "010001101010101011110101110110",
      "011000110001100100110111100101",
      "011101000101110101111000010110",
      "010111010110000101001100110111",
      "001101111101111101011111000111",
      "010010111000001001101001000111",
      "100000001100100000101011011100",
      "011100010111000001001010110110",
      "011101001001111010110111011001",
      "001001000011111000101101000111",
      "000110001011101110110001001011",
      "000111100010010001010100001011",
      "110011001011011111111110111101",
      "100100010100110011001000000110",
      "111010001011001110011101111101",
      "000010001111010011011011100010",
      "010110111000001001110010100000",
      "011000001111110010000010010111",
      "000000111110010111111110111011",
      "101000000011000111101100111110",
      "011101000101011110000011110001",
      "111000101111111101011011100111",
      "111101000111010100011101001011",
      "111111011101000110100101000100",
      "110100101101101000000011110011",
      "110111100001001111111011011111",
      "110000001110011010011000100011",
      "110000101100000000101011000001",
      "000110101001111111000101011100",
      "010100110111000111001101111000",
      "110100101111111101001100110111",
      "001101111100100000100010100000",
      "111000000111110011011101010011",
      "101011011101000101110000101010",
      "100001110011001001001110100101",
      "111010111101000010011001110111",
      "100111000101000110000011100011",
      "111100101011011000000001001101",
      "111111001011111100111101001100",
      "110110001100110001011001111011",
      "011101010101001100101000100100",
      "000100111000011110111000100000"
    ),
    (
      "111010000101000011110100001000",
      "011011100001101011101001000000",
      "101001101111100100011101001001",
      "111111000100101110011001000100",
      "101001101011011010111100111011",
      "100100110100011010110001000100",
      "001010101110100000001000000010",
      "001110000101001100110101110100",
      "001010101010011011100100101111",
      "001001110110100010100001010100",
      "111000000111010010010101111010",
      "000001111001000000001001101001",
      "111011111000010000100011111000",
      "100000011110111101010000100110",
      "100110100100101111011010000010",
      "011001101010011000101001111101",
      "000111001011010110101101000000",
      "110001001101111001101100101000",
      "010011111001010011100100101110",
      "100001110110001011101111001100",
      "111011111101011110011001110011",
      "010101110001111110010001010000",
      "001111000111011010011011100111",
      "110000110000100110110000111110",
      "001000100111011010010011000001",
      "011100110110000100010010000111",
      "000001001100100111110010110111",
      "010011010111001100100111001011",
      "001000010001010011011101001010",
      "011010111010011110011000110111",
      "100001111010000111100101001110",
      "001010001110100100000001011110",
      "010010110101011111000101100111",
      "110100010100110101001100001111",
      "001010010100101111111001001011",
      "000100001011011101100100110000",
      "001100000010000000110100110010",
      "000110001101000011111001100110",
      "000101110100100111100000011001",
      "011110001111010011001111100111",
      "110100001011101011000100110001",
      "110010001001010101011001111110",
      "100101001010100100000000101010",
      "000000110100111010101010101011",
      "001000010100010000111001100111",
      "001000011100001111001011001001",
      "100011001101001111000001111000",
      "001100011110011001011100000110",
      "000001101001101111111011100110",
      "101101001001111110000111000001",
      "101000110011101010100101010000",
      "011111000100101100110011111101",
      "101101100111010011011110101101",
      "000101010011110110110100001001",
      "011010011100001101110000000100",
      "111111001000010100011001101000",
      "010100011100101000010100011101",
      "101100000101101100011111010010",
      "100111011100010100010111010011",
      "101110010000100011011100101110",
      "101010000110001111101110111000",
      "110000010000011101011110000001",
      "001010110110110001001011010010",
      "001001000101000000100010010101",
      "000111011110010111000000100100",
      "101101111001011011001010010111",
      "010001101001111010011101111001",
      "001111110101010001110011010101",
      "011111111011101101110100010001",
      "011000110011101100011001010011",
      "101110110100101111011100111101",
      "001001001101011001111000000110",
      "000111011100010010101010111010",
      "110100000000110011101101101011",
      "100110111000000110000101101001",
      "111110111111001110110110100001",
      "100011010001101111010100000011",
      "110111110001111010110010000000",
      "110011000110111101010010100101",
      "000000111000100000101100001101",
      "001000001001001100010001001111",
      "000001101100000111000101010100",
      "110111010100100010001111010110",
      "111011010100000110001100000111",
      "101011110110100101110101011111",
      "000010011100001010001001100000",
      "011101000110110111110100010011",
      "001010001101000100110101100101",
      "001111000000010010010011100101",
      "111000100011000000000111011100",
      "011101100001110011001111010001",
      "101110001100110011001101000010",
      "000100110011010110010111011010",
      "001000100100111101000101010110",
      "010010001000101100111100000010",
      "001110011001011111001010000001",
      "010000111001110100011010110001",
      "000011000000000101111111100000"
    ),
    (
      "001010111000000011010010111011",
      "111111100011011100001001000001",
      "101000000110011011111010110100",
      "111001000010111010110110000001",
      "101110011000110101111010101101",
      "110010111101110100101110100000",
      "011010000101110001111001100110",
      "010001000010010111010000000111",
      "101100011101100011001011011011",
      "101011101100110111010001011110",
      "010101010100010111100001111010",
      "101110010111000011011010111110",
      "011010101100100100000000111000",
      "010101100011100000111110011111",
      "100001101001011011010010100110",
      "010010010010111001011010111110",
      "001010111111111110110111111011",
      "000001011100010100111111111001",
      "110000011111101101100010010101",
      "110001011001011101010110111010",
      "101000110010000110000110001110",
      "010100011110111000000101000100",
      "011001001110000011101100110101",
      "000110110111101010110000111110",
      "100011101001000011101001010111",
      "010001011001011001010010010010",
      "011001101000111101101000000111",
      "001011111100100110000111000000",
      "001000110111110000000100011000",
      "000110000010101000110111111010",
      "100111100010110100111111011111",
      "000001110111111110111010010011",
      "001010111000010110011110001100",
      "011100110001001100110011111101",
      "100110001000001010000100100111",
      "000010001010011001000111010011",
      "000010100110011000101001100000",
      "000111111111101100110000000100",
      "100101111000111001110110100001",
      "101110001001010011111001110110",
      "000000110111101001000000100010",
      "110011001011011010011100111111",
      "101111001111100011010001010000",
      "011110110111101100011110110010",
      "100000010001110101000110110111",
      "101010111110100000110110100001",
      "110111110110101001001001010100",
      "001100110111011101000010010100",
      "110100111010000011011111000111",
      "000111101000111111001101110111",
      "001001000001101100001010101101",
      "000110010010111010010000000100",
      "111100101110000001100000011101",
      "011110101010011110010111101111",
      "110110010111000101101100011010",
      "001111100111110010011100110010",
      "110001000011100011111100100011",
      "101111010110000010111111001111",
      "001101110001100111100000110100",
      "101010111100010111101110011011",
      "110100101011000110100001011001",
      "001110111101110011011010110001",
      "000001101001101000111110101110",
      "110100100110101100001001000011",
      "110001100010011100000010110001",
      "000100000100110100100000010000",
      "100000001000001010110100111101",
      "110110101001110000111000101110",
      "011101101010100010110001011101",
      "110111001101000011011000111110",
      "000110000000100010010011101101",
      "101010110100010101111001111000",
      "100111100110111010101111000001",
      "110011111111101100111000000101",
      "111111000101001000100100101111",
      "111101011000011000011101110110",
      "101101001011000100001111000000",
      "001001000101100001101011011001",
      "111101110111011110101010100011",
      "111001010000110100100000110101",
      "000110110000111111001010111100",
      "010011111100000010100111110011",
      "111110011100000110000001011110",
      "100010010101100100101001011111",
      "101100000101001111011101101010",
      "101100101001111100111001111000",
      "100111101111001001011101011010",
      "111101010001000101111001110000",
      "110011111100110101011110000111",
      "111001000110001101001010000100",
      "011001110000011110010101001110",
      "101101010110011101001110010010",
      "101110011110000011000111010001",
      "110010010110100001110011111010",
      "111101111110001010011010101000",
      "110001000000110101101101010111",
      "010010000101011101000011010101",
      "010101010100011011000011001100"
    ),
    (
      "100000010000110111111011001111",
      "011101011100101010000001110100",
      "100010010000101101000010010011",
      "101010111110011101110111000001",
      "100101011000001110010100001000",
      "111001001011101010101001000010",
      "100001101001101110111000011001",
      "101010000011011000010100000110",
      "010011010100111110001111100011",
      "111110001110110000011100001111",
      "101000111011011011111101011110",
      "111100101110101000010000001101",
      "010101011110100110101101111010",
      "001000100110111010011110101001",
      "001111110101001100110000000101",
      "011011100111001000010011010111",
      "010001111110110001111111111000",
      "001001100100000100100010000101",
      "110010110100111110110100000101",
      "100100110101111110011111100111",
      "110101010111011001110100000010",
      "111111001001001110111011100010",
      "001100011111100100011100000110",
      "000001000111111111110101000001",
      "100100010101001100101100000000",
      "100111000101100111011111001000",
      "111111010100010110010111100100",
      "101011110101010011110110010100",
      "011010001011100000101101010111",
      "001011000101001010011111110110",
      "111100110001101111100111010111",
      "010100101101010110100110011000",
      "001011011000100110010000000001",
      "101000010110011101110010100010",
      "110011110010011100110110101010",
      "011010111101011001101001001100",
      "010111100110000100000110000000",
      "010110000011111011110100011001",
      "111111010001011111000010100001",
      "010010100110000101110100110101",
      "101111011100011011111011100000",
      "001101001111000101011011000101",
      "100010111110111111111110010001",
      "010001101000110100011000001000",
      "010101111110001010000010000000",
      "111110011001000110110101011101",
      "101000001100100110101110100000",
      "110010100011101000101010100010",
      "100001010010101010011010101111",
      "001111110001110010001101001000",
      "010000010110111110100100111110",
      "001100011001101010001110001100",
      "110111111100011001100011100111",
      "000010000011000100100110111100",
      "111011101100011111111100110100",
      "000011100111110000101000010011",
      "011111101010101000011001111010",
      "010010000001100001001111010000",
      "111111101100111110011010101010",
      "111001000010000110001000111101",
      "101110110100011110100101001110",
      "111101011110110101001010100100",
      "011101110000101011001000100111",
      "100110011010001111000001100100",
      "010001110101000011000111111010",
      "110111011100111010100100010110",
      "010100000101001110100010010011",
      "100101110111111110111001100001",
      "011110011110000000101011000010",
      "010010000111101111101001001001",
      "010000110110010111111110100010",
      "010011011001101100111100001011",
      "101000101001111010010100101001",
      "001100111101101010010101001111",
      "011010101000100011011001101010",
      "011101111100011000010101010000",
      "110101011010000101010110010101",
      "011011101000000011000101000001",
      "100010111111111101100111101110",
      "011000000010001110110010100010",
      "010101100000111000011110111011",
      "101101010010111111100000101111",
      "101100000110111011111011011110",
      "101100111010101111010010101110",
      "001100001001111101100100001010",
      "001110001011101010001101011011",
      "111010111011100001101000100100",
      "110000100111101000111011011011",
      "101011010010100010111001011101",
      "110100100010100100111100011100",
      "101001110111001101001100000010",
      "011111111111101100001101111111",
      "110000110110111001011111100011",
      "001011000010101001110010110111",
      "001110011110000011111011011100",
      "011100110001010100110100111010",
      "001000110100011101010101001001",
      "110011010101110000011010111010"
    ),
    (
      "111010000010000110111000100110",
      "000110000101100001101111101100",
      "101011010010011110111100010010",
      "001001010011010010110001111010",
      "101000011110111100101001110100",
      "101011111110011100111100001010",
      "100010011011110000011010001111",
      "010010101110001011011001001010",
      "000010110111111001110010111011",
      "101101001001111111001100000011",
      "010000101011010101001100010001",
      "110101110001110101100000011101",
      "010100100010010101011000101100",
      "100000011111000100001111000111",
      "111001111001110100000111100101",
      "100000100110110101101001011100",
      "100110001010101100010101000110",
      "110000101110011110001001010010",
      "000101001011001110100110001110",
      "100100100110110111101011011001",
      "110110010000011000100111001001",
      "000111100011011101000100000010",
      "101100100011110100110000001010",
      "000111111001110010100011100110",
      "101000010111010001011011001000",
      "100011101001110101000101010110",
      "110001011111110101111011100101",
      "110101100000110101010010100111",
      "111000010011001101100010100010",
      "001011011101100001010110110111",
      "101010010111010100000101101010",
      "101000010000001100101010001011",
      "101010101000010001110100100111",
      "010101110111001010110110101111",
      "100110110110010111110011001101",
      "000001111111101010001000010010",
      "011110100110011111010101000100",
      "001000111111110110000110010001",
      "010010100000100000100001000000",
      "101000010100111110101000000000",
      "010101000000001101011000110010",
      "000011000101011111011101001100",
      "010111001101110000000110111110",
      "011001110110101100111010111101",
      "110111000100111000000100101011",
      "100100100000100101011001000000",
      "101101000110111101101000100011",
      "101100100110101100101100100000",
      "101000110101001110111011101011",
      "100010000010010001011011101100",
      "101101110011110101010001100000",
      "110000100111100010100100110111",
      "101110011101001110101111011010",
      "001000111000101010111110100000",
      "011101011100111101000111110000",
      "011111010110000011101011011110",
      "010011001110101010010010111000",
      "000001000100111011100100110011",
      "000101011101111101010011111011",
      "000010101011111011000010010001",
      "011010100101011110010011010110",
      "100110100101000100101001101010",
      "111011100101110100101011110010",
      "011001111001110100010101010111",
      "110011000110110101000100000111",
      "010011001000110000011011100111",
      "111101110010010101101000100010",
      "110011101000110011000000100110",
      "110110011001100100110101110101",
      "011110000011111100000101100101",
      "111111000100110000110111101001",
      "010111110110110000101000101011",
      "111111110000010101111001001111",
      "010011000011010011000011011011",
      "011111111011100010010010011101",
      "101101110001001100010111110000",
      "100111010001010010110000101100",
      "011001100000110111011111100100",
      "000001001110000010011111111101",
      "110111000100101011111101011110",
      "001010101101000110010011111011",
      "111011111110000011001001101001",
      "110110010010100010001101110101",
      "001111011110011010110101101011",
      "111001001101010100000101001100",
      "011110110110011011101010100001",
      "011000001001111110001000111101",
      "111100110011001111001101011000",
      "111010010010000110101100101010",
      "111110111000100000110110101000",
      "010111011110111110100111100110",
      "110010001110110100101100010000",
      "010011001010000001100100100010",
      "101100111101001111110000101111",
      "001111011010000111010111000000",
      "101111100111000111011010001000",
      "100001111011101000000111111000",
      "110101001101110000111001001000"
    )
  );

-------------------------------------------------------------------------------

  -- constants for State permutation for RMATRIX
  type INT_ARRAY is array(integer range <>) of integer;
  type R_C_ARRAY is array(0 to 3) of integer;
  type R_ARRAY is array(0 to R - 2) of R_C_ARRAY;

  -- number of columns to swap per matrix
  constant R_CC : INT_ARRAY(0 to R - 2) := (
    4,
    3,
    1,
    1,
    0,
    4,
    0,
    1,
    0,
    1,
    0,
    0,
    1,
    0,
    1,
    0,
    1,
    0,
    3
  );

  -- columns to swap per matrix
  constant R_C : R_ARRAY := (
    (
      94, 97, 99, 100
    ),
    (
      96, 97, 98, 0
    ),
    (
      97, 0, 0, 0
    ),
    (
      95, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      94, 98, 99, 100
    ),
    (
      0, 0, 0, 0
    ),
    (
      97, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      94, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      97, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      97, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      97, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      95, 96, 98, 0
    )
  );

end lowmc_pkg;
