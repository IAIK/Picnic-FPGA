library ieee;
use ieee.std_logic_1164.all;

library work;

package lowmc_pkg is
  constant N : integer := 256;
  constant K : integer := 256;
  constant M : integer := 10;
  constant R : integer := 38;
  constant S : integer := 30;

  type T_NK_MATRIX is array(0 to N - 1) of std_logic_vector(K - 1 downto 0);
  type T_NN_MATRIX is array(0 to N - 1) of std_logic_vector(N - 1 downto 0);
  type T_SK_MATRIX is array(0 to S - 1) of std_logic_vector(K - 1 downto 0);
  type T_SN_MATRIX is array(0 to S - 1) of std_logic_vector(N - 1 downto 0);
  type T_NSS_MATRIX is array(0 to (N - S) - 1) of std_logic_vector(S - 1 downto 0);
  type T_RS_MATRIX is array(0 to R - 1) of std_logic_vector(S - 1 downto 0);

  type T_KMATRIX is array (0 to R - 1) of T_SK_MATRIX;
  type T_ZMATRIX is array (0 to R - 2) of T_SN_MATRIX;
  type T_RMATRIX is array (0 to R - 2) of T_NSS_MATRIX;
  type T_LMATRIX is array(0 to R - 1) of T_NN_MATRIX;

  constant K0 : T_NK_MATRIX := (
      x"c24f16269830180b15c295c21894889c5a4993bb70b1c39f0237d95c1e832002",
      x"f640e924b648d06edea78046da1e78a26d71fa9440860faa4cbc257c47d3c096",
      x"3d3695b840d6075fceb9a455d71b25de18836fcc47d605fb1fac80409daf26e2",
      x"8a271257d44205a985ded37c470836d74ad0e971324e3b862a3963a5b9c4f7a2",
      x"df2eb407ce27572ae41fdcf686bc11d061599c6db147d4e978eb04804e15ac95",
      x"b0e074126637510f3107c01c2c656372546dabdd57d3cdded8de215d348956e1",
      x"77cc10270234b8eab976eb6a7bc14c9e73a12c6b146c71f3aac76cd76f8df8c0",
      x"7bbe18d775183d8345ab2f90bc3dd0febc5bdd2860af20aa44ac6b22d5c5e32a",
      x"830d1ab541a7d07a3d98adf8bc3e15b30a9eb112e2ed341593fa95cc8f83a049",
      x"5d25139cdae197e627e4d26db6d50ae2294a8e9ce384d6e3f20965fb2edcce00",
      x"7238e686f74aa3d30d735a6e88d501686e8a54c7583996b20e7115685cb51cbd",
      x"5ddd8ba2053277a1c6360cf4db4378c956836e9514d0d9c3451432a14df86dc7",
      x"3a2d05e8546d93c5e3ce20a26c95dfab010a1abe69d22566badbeda186132eff",
      x"2b0ce15778fb6c90ad140434ce367aead4c659e347822d26275dc92cc3a616ae",
      x"423824b58072d20426cc26bec22f1f3a5465454a7e864bdbe19261b5c27e5cb6",
      x"db065668b86a73d41197250e1f667ad3447db4b113525e0375cfdfc9471b94e2",
      x"f9531a29cee0291d83b2cfbee6e9306e099ecd3146796c28bd8cd97803eb156e",
      x"a34178670211bf883a60223864b86dd9294a14840a9ab08a3ac4a1f44847bc55",
      x"38a8892657bb861c65257754b87b9d297b41b2db0d8ed147cf7e8a958e5ecbf9",
      x"25495e9beb966e72e83880922fb678c2ff91e581b563f9f2b16516321e12a707",
      x"584c3e22cbee4b51cfcfa8902c657904f1b0f6e9f37ec763f890e30e3f238d4a",
      x"8e5b76495103200a6c606607fd4842ebf5f2c826474028e9af9b169ef27cf5f2",
      x"45c2b9cab066791dc533a34ec635f438f7627c146e04430918ee12333ce27718",
      x"dd6d8a359b033f33053da7878b7ae6bf0d340ca47bd549c94313f318ef671179",
      x"1886654059c80e73cdbd9477835c0f9a069b6a323fce5ed7a771d981f4080073",
      x"ac58c02e866ebc9abb0af12c99a746bf35a0b342bb5648679cb4076055c83fb8",
      x"4812a840b13151f53d93641d7c300fd1219be4b8cee9a5fb115fc08f623cd847",
      x"15de9bf62f74f7844f39b049712a8f88d7064f2c8cf6f4252b4b31564e352705",
      x"697b604cc8678b12f3394e0ec80120e2efb8242270ab8ea7c2af2ba5046add11",
      x"42b1ef0166f22fb094bdc91abd6b6a1bb56aaaf6d440ffade3dd959ff43c6139",
      x"2f7b1dc3d1f522b03b1bba8d093cd4634459162ca9d1b571feb93419fb3ee9ff",
      x"9c60f72528fedcba9213efa8eab9c3f9427ead5bb95afeaf50aefca690790061",
      x"00996f849641a73e29292a1cb01d0e9426cd1ec0167a4bd1e93348f0deb0bf19",
      x"499b674e47658d70a9ef34bcc5eff568c4518440ef0c38dd1044bf14bf529b58",
      x"3a261a45f9a2629ed52f5c5060c2ae87a7929ee4bd8cc177b0d78f7d50e159af",
      x"240edfddaa2cea8e4466ce493fccff26b3a60c883e7a3896becb9df8e77584e3",
      x"4404dc19db5f5650f18fd0f2164e899c27a7acea565184aef342742025c05df6",
      x"a460f29d89f60a5bbfee3ddfd1b6e62bea592421d0a14c5418b1ef9e0483e777",
      x"09c1fe7d3c232251481d0762aed68c9d9d2125a96564b258c6e087289c9e533c",
      x"7eb54d97df60a20ec4efe0f90c2e482610063630efdb6538a965f6603598b223",
      x"a7e14f3e7eb11b403e3d91d4d5c3fcf66282a4861d628ecf089e942b09954e17",
      x"d5a6234032fecc09da57f7c288a0ff2beeb267dfbb6869b21a757771d71eda7b",
      x"261ba5c44ec3ea425391146e389041b221dc68a2ae13eb1124ef34a18c3bd9f9",
      x"5aa5ba5ce9fb227c597e4ed12f13439a66ffaa10876d90967083e6f3d77dfb35",
      x"f1702c44ba077301d88a8a30776e2d4b26bd61a6588343c936cc0b6a116ab01e",
      x"dbadcc7268a212e12a46fee16d4abd86e08fb1265634edb47d7ff6b9597c80d0",
      x"01b9615abf0c900b78ee086c8247ac98f70227697e50463e085b5c8117efd76b",
      x"5672aa4ba762631a073850d035f03c7958d7de79f716d00edfedc4bad6d83d8e",
      x"e2eb32a1779adbb71ab641c076b3699f2c672237cbd5e673ab97346eceedb5ca",
      x"ea77abddb3ab8d1b79226840ea7ffafa4a2a12a2bed46affd8d3ed5383d37cb4",
      x"aae004edcaeff2df5a4d5f7537a89f7f0c6393a7a3f4056e9f71a869d47b6da6",
      x"2f6a4a14d675af4f62a09bcddfdb7310fac2a45514263a9196ef2e1854eb0f78",
      x"354ed7d5f3c33d10c4037386ce9acd68029be252861c6a2e0b2299bbb83258ef",
      x"31dcb6b20f2731df54362af0ee3f8064e0f4da0bcadc1fbec7c6cbf539dd3894",
      x"2a76fd866e09fbc9802ce6753064b3086cc9aa7ce7d93b007f2fe87f95927906",
      x"57fe468d84b1c0a65029eec408111da95b33bf49c99a4ae8b8c7f27575194766",
      x"13d58147848e05bfba9f5fea9df07061dc50003ff6ea21423ccd4d87146a531a",
      x"810f93c83ce59864cace66afbe4cf9159198d84c55e458d2cbe42f6317b104e0",
      x"981346e4523967f263748511de88dc0c9b09a344f7c9a12569c61abec116cc55",
      x"fc5c2cb25e5539545f97190c85d0e66bcc431aaa731e7e46226736a500ebf79d",
      x"7cb624cc7abc85c94928e9b55c764936b208a64b8c242d82c509fbb8e2044bb9",
      x"b25e824f997116505ecaa3fd2f3bd9af81f463e9e013b897903810872a5fff17",
      x"904ef3b39d9cf163e470978508d8cacb6bd6ec395aec35f701ebb9a6c266d4bf",
      x"237985390713a7dabb4a1a33cf5ec359c5c2befa603b51ba818bcf1a00d2dc43",
      x"14392f4a50527346edbd3a666245d64619a5893e1c569d1f97293a1557d6e835",
      x"fd7ef5fb9d113f8c100f12d0ca596f8a916e16115fccf32b670c268dfa5ddea8",
      x"036a19bff4ac95b845d4812836899e1919acd429fdb38b0059673e4b33c8aa62",
      x"11a74e863851a986d32f334196d67819d34437eef1103b48c1a42116752e1f5e",
      x"f7117fcc9d5870136a939ce76c0886c5c315447808cdf6704ca90abeec77d6f7",
      x"dfe2b8fe2524c95a2444597b96bf3c304fb35d20d14d7288c5ac19d57e6e3809",
      x"4dc18c6aa69a90106a8de8827ecdd9783247ae8b6a68aeb56df09e4c57cb1713",
      x"2c3197916fdee6480393ddfdc9786756819099bc0f14f02c6080245e9c81ac8b",
      x"8fa1d9857a8b1c9a97c29f03af6c8e48be8c8e31f206b2a6bafe921af83bd522",
      x"40024e38234de27d7186edb79e0d15ee96050e0b4dbff8faeb3dd93def86b649",
      x"5f5ddbab5d343a445b111ff0aec77f137cae6003e97b16f39f22fa90267b56bb",
      x"d6a0a3bed34676abea4bfe3e575fbabe0d45141f50b2e2577c86a8c3377280fe",
      x"215bc47fbba2de00b78c0d6a655579fd08214a9b0bcf39040d1cc5cd25640a06",
      x"1d1d439947c5518111299d4cc45aed3d2850df28c5361f774e7fdc4550a312b7",
      x"687fdf52ad40235560450a0789abf5480c21f6fd5dc544664e302bff6db81592",
      x"d2a187ea1cfce06074d796ffb9ece0b71895009824cd9076bb752ce8c75a076a",
      x"8825007263782bfa7761e87bab61f5a4fa5532a4f464f2db6fc406d30c7fe15b",
      x"79a1105ff7cf0125f6c9b44165afea7572d6348a73697937d8c400a5985a6a54",
      x"86dd9a95675cb82a557c3806de4e048c218c2d43d1d6276ac462890d70c7dba6",
      x"2fdd71ba44fa4caba99ba6b4dc9794ccbbd0fa951a38c3465b8dc34115782072",
      x"41a6767be5fbafd83fc5f0bafbb4d7025b82875746bf9596aabc6a6e572cb39d",
      x"b406cd54971d48fda82b563b89ce6b50cfbb9ca77c7444946f452d9139b1b59e",
      x"d6ef21482156f6a2b361983bf26d41359288c03aab308fbf9a7a34aeb4407715",
      x"8986be8ee9b8f36adf3012aa2a619ecde57e9f1e11781ed3a1e2a1a3a9b1195b",
      x"b39d58f9fc03ae17e8c785dbf6555633f92d8fb932450c4cd7060568c003cfb7",
      x"f931c22e85f8a9a2a76fbd30d4f50adb0b9dddd2d8997716512dab8314277489",
      x"da3960fdc36656482786206945529d4be95f900aa1919a483cbdf9c7d0cf0ce9",
      x"b92c60e94886121c4b2d219bf904fae5ea06df7b793e5498ea8836aa8c743a9f",
      x"18051b67ec7a55f9587bf6f82685865c9bf847d60964351e255a79ba57e88fd7",
      x"c99d0eff7bc04f823e874d02eb475fc8cd98cdc520354c89b3bc206c91a1f4bf",
      x"95a2b0c6872c24418a01f2f05a76f0a7023064d492bef254f7194734c32d5dde",
      x"6a8977cc399eb408cdf6c9540079a9ee3f12151b43983fb3c9d382fdc27f2a27",
      x"c33fcef9c4fbe2c5902393a5eff6a8aa67e1111d9d7db4b3d4a64d02f8335762",
      x"c1776520ec7fc37142faea44c71cf248d1c74679db32dad31152400cd8f25de2",
      x"ed80fbbb08fc7e300933e609ba903fb8fad082c26b843002446344e0619b3175",
      x"6afcab88892f7b6eda5c25959c854194b20d0186f92b199bf29a574b308f23b4",
      x"1b02bbb0be7a9a9bc175c99b5b02020263bbea84937f5e91a597c5b1ece784b7",
      x"4e567d7b4524bef27ad261a20e81dff535ba83fa742931c9f726287b5615651b",
      x"0a60bfcdfd7430d1a4cb2908ef44a7feef1d0bdcb208c4c9a3f624910edc72a6",
      x"16472baf01170d8dfb16f57b45baaae5dab527117bceee32205b0217034985ef",
      x"cfb2e3b9c99512eb00e119adfdd771e6fc115a172ff564278f40186b51d5fd7e",
      x"1a8b06d4283d3ef90bb8f04afadbfdf2e4bbe44695ac0a53056abbbebf2d24c7",
      x"a513d6803f7a04e20571328d3b5ee408c82fc8ad591559beb69d9be896aa366c",
      x"cb97035fac89616207c8f233abc7f794b6fd42daed950757f5ac5d2ca303e639",
      x"7ead7eb42d46bd736b58f8111fbc1eac0f91927428ad7762d19882462aedf8da",
      x"4851a50a01aaf0ea1cbb9c945cca53b2718556fe687429246ba9a77facfacb8b",
      x"5af275ea6784361d60dc75a193388cde3a94341d26f32bec6983b69a4dae2f02",
      x"f4ea5fa9331581f449a9c4cdd53294ecc16f0dd5a76b75638fb9822d1ba46e18",
      x"1e7863a3418177e1a5a9ed0603da0052a70f87e5f538000e0d922ab1f1561021",
      x"69749ec04081b70e5dc266eac40a63129f857e0df2e151c673d78181e3effdb0",
      x"b05a2216f3f75d2b5e3a9948e986dd02af169c7c8319f5aba7d2730c57a6c42a",
      x"9374f0d5dfc7f2ea68398fd7120352a1f8ec1880e21f7d95cd6abf4f332cbc8f",
      x"f798067862521b33d3fc02c9ada8a59f921460b683bf4f556775a20380578277",
      x"b221a29a9314a702b486f4ab0e84467712c718751f54b9914767521e66893fcd",
      x"5bb9e8c44619ee4ace310e7d9366c7da3c6c379e66aba1eb1077df989d28bbc7",
      x"02f32ce2a965d5d3a2485d4291149c20ad89963bf385d5bbde05eec91de522fe",
      x"73d78621ff81f8f40dfc9d58c6b2477b8d99de5077eb7372cc4a043273128b7f",
      x"397e122c24e7ee52347eedbd4eb9a092c9c9da9414e75150f2e22fee644944d5",
      x"fc1e2a5d8a031d87112efa103e085ddb2c2b82ef283a8bad49a98c0da754e1e9",
      x"7db391a39f125e896a009de0993cbad264a10f3828fa435bd68ad9baee084bb9",
      x"b9c0bbb4e0833e86fa98888d671808c831bb3769a8b1c8fe6ddb0d19db4c178c",
      x"d0d7d5b15f70155070dccdab5574ddac32eed2284588f399c07b5d8ae53ed7f8",
      x"8f4d9cf63227e9bdf3614654665a218f90f011268a0ce93013720dbed8b14f1d",
      x"f32f97e57618f37bb06ec58d91a9b2e5d08629894ac29c56efbed08598a17094",
      x"3a887024e9a4b7dcff9c541d3f843fbdd0b2f4797c32be2f197507abba16b2a6",
      x"c3b0343736d4135fb53553886ae1458d3fd85aa66bdc59149dfa5bea1345b488",
      x"7a5da86422f8d4a15d372a745840f2f638d909e971b27a8696a6e51529eb2523",
      x"f2457cc62deb7acb9c7abb580866c3dde0c47365ecda84599b8a509887fc259b",
      x"7820e0922b70be17270c4d2b083ffa4c8d0e57da0dc039af3a7d540ff8aa69a2",
      x"1192c123b009c30c53a9dda7010bf753307d7dc3824c9ae7b2f8c8949b622bb5",
      x"55a9298805c6d11f09dbc93265a834c1bd082ab38ec9091898d38670179bf691",
      x"2b5635de5af11a5419333a66ce04123024e1ede6298781f7038ad138bdad7331",
      x"b6491aded1c367411b77e215fa87bcfbd47f70e31fb4c8032718810b4dc4d969",
      x"aa4eaf7e6d91ae8a196b9b2f52235e15e9a0eaf966f78b5d2f3b2c1f4cdda34b",
      x"73ede0474e1cbdf031993dc9968e237dc67735a9796cd9df0887e4b1be62333f",
      x"9a3d9abf51a2ef22fad113bc324c5d8c68d433868625e3cf232a01c974f60327",
      x"fdf0e00d410437fb60ea23aed0719dd3cbbab32c0103b45a51fbf267d5c759b8",
      x"e8f0f9065b84913a0da5fc9357e830ac4c7328fe825678a639fb9442fb5766ae",
      x"e930023fe1daa33e0178b1b11daaf6cbe9442249811a61a2c8802fd555f98c5a",
      x"1d1c8a5e9a239044acf85f61124debbf190c5c6a85f5dc7ba7a9b255c53d7af4",
      x"0d53672941a259667661819cf575fdca47b374da46e0d7fd4ae8d3a364233b30",
      x"53612ef915b99a475819bac78b2e15e17d94156fb11e54d446af642835b0d142",
      x"05f766119d68736dc037876adec0d42217b7d57a9fc8cfea1b173cea0e1351b3",
      x"891f9d3ce4388f78be186fb978cffb36c14645483e38fa8c003e3d43ffdbd52f",
      x"bb9700d98d6dd7a1501b99f2fd9e4f77a44d52a2ebb73d55a49d1ce5c342cc53",
      x"59d7430f9907d890a6b0e805f34e54dcf7c84065a6a0c02a51663b3f7abf2ef2",
      x"8e3e1f6f83c508b206ca21c0644fb16c032544af4210489cf9a58e53bb4f1e8f",
      x"b571c3d7aae35cd8b287392398afdee8ce3234aa2dea3785b5c390df7d2ca2f3",
      x"02a3d32a6af929d2798573591c927b0bf7c127f7ba43da82179668aa079f266e",
      x"416cddd788e30712f02f34783bd97ca90625d1f47aa5c177c681135e09baccdd",
      x"0b563c9b145cbb236f8620bff80742c4c95af31b8848cb46679acb1b91df6b0d",
      x"0ef48935e45d6c5625bcef9f856eb75b2414bd1b4a86a4b9b5169fb249a528a3",
      x"85c0e9c19bfa2f798b6aeffd9d84ebde1a702003a47a8358460e66e3ce000b02",
      x"8db02adbaa1a1a0640ae43e27b368b3250152680de465b9824bb0f6a698cd0f4",
      x"aa68811258eff86bdaaef5aa996c32e1bb59378c19b655222a50dadb3723fd3c",
      x"f14b75b894f34184e420cf9ce0a2500caffabc1b4a98046f5517050c4cc2dcfb",
      x"e7aeed11ffc83a73ba2228caad8e3cdbbd0159deff414ecc180bc62e505aa192",
      x"612ff3dcd8082ef959162f1122dd9e38bf30537147372255dab4c34e694b32dc",
      x"9ca7bd869c86b680ea9c9a83979d07ba8dc952367704282a704cc4466b920f88",
      x"6317563cd43e1d50aabc1b48c9d08d1d59bb32c2dbdb2808a107a45acaee1ee3",
      x"10cbbe8f9b6a8e30adb7df4da7301b209633c012b5f6b39471457adc7da798d6",
      x"1e18062aaeee9869634cbdb093ea3f5c6300ef8bc9d29e740c825bb59bea3275",
      x"0a90ae9100d543ee27fc3d77ff2592ae0cd15b96f4a0e953adde812229f9b0cc",
      x"682b5f46ed5783fa279ffaefd8c4978b525d38b6fd0dd92c78fc03cf435bff9e",
      x"f98fbd60b29ad3e3484156622311ba204e74af280ec2980f5d0dd92660cae053",
      x"497ffbb2851a519f5205476cd66197fdd68411e07f0360b70d10556cd8861dc5",
      x"21ff31b077973ed991643c4a1adcef23cb4f82ef91765b800f19de4b70df271c",
      x"1968d76ab25a642c559976eab4ea2c8536dc4ab1bd2d01d19b0368224ab42845",
      x"6f6bf4a6c66b70989578919bde8a2b3402f2a63139806fb9cce8a19f69de11f3",
      x"a83cb1b7e0db0300ac5bce11818b7ef1cd89bbda3ab9bf14d3ce8848a178b734",
      x"ed1a7dc8531ad1478cd0769933ddb0d07d773b47dead0236696f01b3d423fd04",
      x"60d45bc3827bb368e28fdc8e56773d948ec61d5a54a69dd2847cc03b51e0cfa9",
      x"90ed22afd844307273a42a487bb9497600da6476eb6715023722dc270b3e8c89",
      x"30af9ccfae1baf7347c687151e56396718a3d5433e18f62e22e4e0f46b05e8cb",
      x"88589764b906e8711fc33f2fdca975955a16d97fc42273a403a4e9ecc5af034b",
      x"ea3b2360ea309af860fe01a91d94cf60d7b595eef010787acba17046693af597",
      x"1f520052f729e1e63479b23d65c8dbd68ac90f703c3f25dc0e69915e18749925",
      x"b4095731746c79257502f447988786a6441db0a33891363bee73c5eafe0b9b0c",
      x"81ee3a3c51747f27bd57c78b166d5836571435b4ed26e5563bd4af441cec5b1c",
      x"21e6b299ae8ae1fbc0ac7d65652987809759c10ccf22bdf2041b25264d26e5c4",
      x"55544f0b1dbebfc798614bc84480324f77081b1007b704f510f2508613399864",
      x"fe1e600576be6ab4a38bc12c11f33645c569f565cca8165562aa1e685a5034a9",
      x"c948e24859380182a0660c011b136f357ef7b5355b105790bcc03b351676b7e1",
      x"b1f8fdcf882e6737597768cd3c85dd300804a28c232bd6c2033cbef43c3691b7",
      x"6ed5476bf67de705c7658c03b36b9b73ebd70964ae402dbcfbd778adc54ed522",
      x"2e3c1a05ec74e0a6346622b271fa23b2ebb924da07162cfffb8293143edc18c5",
      x"371fd3e089b3e4c9c1bf8a63c210b34324c32a53832e0edb4cc2348882b2c528",
      x"4fb1cf41d41839e19b0c7dd319ef6e3fc31f1fbda9715a76a85365337f10b7f4",
      x"cf14bcbb11aa1461ab2be4ec8f79402268d396b9e3471bc6e3880aafb43de84a",
      x"0ccc9af4226cf85296d0e7bd0a6c2039599bc18a62af614e55cc7e01e322d889",
      x"0265145a29d67c7fcf0af861abf41a15a544f53059b5378db93a5cdfd2e75ec0",
      x"7e280d145f7e0f457eef7188d8cbc4250f6e3043a26e33a43be142152a5a280c",
      x"b80433b672cd5e577c1c2a02f1b5fba503d01eb19ac8710b15faba8acdf15a4b",
      x"c0a93db2547f6e534f6cf781ad1fcadb08b4c1152ae4f9a22e78561200aaa927",
      x"14748261eee7ff017134cc5389ef2977eb08deec1e4cd69b0bdd5785fabc058e",
      x"2188f184443335d6a4a51da7e57d4a6509ac7dfda5e3587568bf1a04bf81a01e",
      x"b0a9a7018afe39ebcb8875b17bc5d6b6b275631a1a5f4aa14b4ec594c2779fbb",
      x"27df7ee4b33454b92a81288c9e8179c6f5115efa03e0c1f6f36809cf5e00a5ea",
      x"f619ff5552bddc2d55d1bad6c1ee55ba01d47e6f81c1d1f46c4c8a360aacb607",
      x"20c220576216d59f8eb24d35c0d6f514bfb9a0ad5971bba5844b73dcb2dad27f",
      x"4f91abf8b1d2caa484e6c3f017c80e31eff8d6c5f0aada36cd4320620cab5eb1",
      x"748b8bafee6816e5c300bec8ce520aa020ee356db7c444ddb6365ed5307e4f1d",
      x"67f5aa3dde1d55d4fee429f8ea65da2ee776ec10a1aa4bb454e019b50e4106c0",
      x"83793c6f8fe863c9d6af6b8df00fb51d22c446fa6b22445cd98453de310bbc80",
      x"0dd3fe2cb900394dfaabd69413571f2d530378b902053f48c44a91343ef8190f",
      x"3848be5eaaa50f757015426da48a5dfc97c45f152f3acda387db7ebe57efcc50",
      x"7cf59e00ac657f48b5ea977460381431d00f3e3f42465fa6acd09f47f9301f3d",
      x"3cac4d3677766c3a73b307ca04e9343f298a8d8da431f2599260f2c83305a0c7",
      x"2a530bc5268afc39cfdb268449ba81978b8085a3c0a7d89f9a7f69d6c4f7fa8c",
      x"6e7b7d387da6f9b85bdeb0fb2a267de333d8dc4c7d45d7ef63292a4407d9db67",
      x"f592e0b756db102603fe4b1158afecb88ffa23ceebc4e04c18b3fe0401ae4809",
      x"b5d6b44e4485ada30c79e7a6942f3ca3fc85e2cb97bedd32496f2d1c5e1d3adb",
      x"edb9ad325dd1294606a4bf236d6c1d1e762866ea870114da595ec331b4da66a0",
      x"3ef09f7f572a348a4fc5916859f24fd12abee5ef05430c985e9f87cb222cf274",
      x"7f5595b2a54c9fcbc06b999d15e443c00566259eda7ae241473730c04ef71134",
      x"70bd2db718c426b22cfec5f457ee101917d246eca7bfe8d607b1f4258d36a242",
      x"3afc6f323afe007f6cdb08591b618d35fadfeb751ecef77417504fc12d4fb065",
      x"60d774100b0b6120d0af542b712321ca79f536b33d3174a8af66d0e951d93f22",
      x"b134bfc37994aa37694256fbdb3e5f6131963e3a39f459835c1a92cff40b9182",
      x"7ea409b8c4f2eb0e927153d2d8eb016aee9f674db7cb2b3091c9de7eb3f4ffc8",
      x"10c53323d95f640a01a3d82698101792797df02048fc40ffd3e75f1c489aec3b",
      x"b2813c320d1317fd795de01786962f75781584b8c46f69980dd60740d6a1d5a3",
      x"2cdf292a2ca16fa501c12120c4c7d11c337e627681980a65ad53f7eb07eba3f1",
      x"28b5fdeaf4eb321b06652b6af6cdab75f5ea7adf452dbe0a65999fa4963eda4a",
      x"e82e9ea869dc5b16f09bd78d32cdd7affbabd8e448c0045546a307c9650de301",
      x"9f238fe626397a49d29ba7e7af74052dde05d1c41dd2169053e2641ffc261134",
      x"3a63a631ca5f6c2a6d682a9d56b7020f9b68a000808030353acb390633b11ca8",
      x"46c2af8646670d4aaea1172c2506bab0539ca844ffa0d694a1d275c4e32db653",
      x"467f350eb7c6071e1b9a4b430d5a45027be9626b0c4d26ff117ccb48101fb522",
      x"608c31ee9bdfdb69196997ee83de9687189310587870d8338aae7ca995762c01",
      x"fc300b3ade38206c2e1d89c35486e77504a7902f6d0ef1a2712a1a393c86c79a",
      x"61cc38aa1bc9769b715be42a2869eea41f633a94dda743ed75a0787e388f1903",
      x"751725c00de65176462c2ada99649149d17ac4ed6944b7f083376e8349a4b02d",
      x"c24f8a973fde4e125ac334ada68fce7ff3c2ae621dcf36c9e89428eaf4f5f5f4",
      x"218ee9bd65ca84c523d6a0543a2fb0bfa7faa151cd07a30c6b27feec289372bf",
      x"f300c8f7d097ab163250e4aea55bc3da6f3a1ad7ea031534210000728c071539",
      x"c7d041ce78fd6f902847590ddcf3439be05dcf030b3227a2375c2e12da698e09",
      x"c18f081782e2dd58db4d70f7bfa06a815e7eb1a73a85f258ad884e15f33fc1ce",
      x"2121cb6a132c89b34f26f6cf0e9d4de05da4185acbdf55e55cf0b7c02ea3ea16",
      x"0068847ad4e991602d4419c55399098671c97adbad79d44c2928b4ea92eff2bc",
      x"f3e1b26912955775176c54f2b88d002d01c71d1d48df40a8c8c6ec34f2b83813",
      x"ea8e94fe55a837e33a6a48bbe875eb0091c01e0658976b2901f525a28101ebaa",
      x"45d61c762b9069022caf77f7722210ad0863f4a7757d2827da066c3ef6dd04b7",
      x"51d8c014a4fecf76a3f61edf613000e55f19686d2e0c60406de91036af40c2a4",
      x"b391d427e0e3b2cd9d47e0995f88757644194288490dad09a2fd3531629de2dc",
      x"beeb8c3ec4eb66e359b090c834ba0405be2ff0e13bb62d989ce513b9f033e007",
      x"d9c12f04c69c0e4a38f64cd155a946a1673e6f0a6f4a30190c8a933040e9ad0f",
      x"e30423d54628baca33a2218432e3254757f3e316ee4e2bd162af696eadaa2493",
      x"1659ee274a9804f1b7eff750bd8c7ebe3315a3f9bcd697195db116d6987fb120",
      x"bc370d915607acc8ae95fa3eb9c00a1896b04e934b96f2cc36b6729bc5586bc5",
      x"402ec45dd90fba346d46fa5c39f4dd819c05db699719e231332bd4607aae2e8f",
      x"7b20ee4a112b9010d2f27f1989852776b5732ad7467d849073f4e6e922b36731"
  );

  constant KMATRIX : T_KMATRIX := (
    (
      x"0d2f5f5f3cfd4463eb86738295cd0f84b4da42a6db04bed6913a373429b9ecee",
      x"c720f317af787853b1d1f0ea110aef330acae297d7c5855f40ccd73cbdb80e3d",
      x"6f789b4e07eb3dff4fd4a902de924ced9aa618554deaf8035e9ab97e660ce1ce",
      x"ebb36404920a76fefbd944f2a63aa33ae2558c807dcc29ca5ce706247c23f070",
      x"cec02aa03a4390fc2bf7c0e5fc2be3d5e73a819bd064a170a1d102206b6e0c4c",
      x"c4fe705a6418e9dfe445736e903c02a6a364d881d9914cf4cd8393852a65f04a",
      x"923481d4ea338f64693065ee03f652511578ea9f0b17e1ebebc5d552b861e2d4",
      x"253531ab5710882a2867589d5fa3ddf9db951ce524cbd3a9bbe590c4663191b4",
      x"b806ae845f30a73d587665a3cb4460955d01489e4face459ccc291f37520b809",
      x"e3666b84ee7f1caae7d57016465dc8521747782b32bc5806f9d8541b3ef3d89f",
      x"ed78860c94c8f156805697154988a021a16a3a86846df7971af85b2bea7e6460",
      x"f5f0aaaf3a9bd6ca7be4d1bcd0e4a64a0e5e30751d5c7f4804b540ab07dedffc",
      x"00c3d99b4378e6c39292feebcf58e772d31f6526642e5a2be079a3797ea4a25a",
      x"10990154edf80eba34a416a0f5d6503cbd85ca2168c2d9fa7baea7682e6d0d33",
      x"aaa67a26a2c81501abbde83f1b5d941b245af57e96637bbe2a6c2fa097f86eab",
      x"5f27de53b4c30557bc9f0c833f1466938445ac4dfa5cb52e28b26de77b80e6bf",
      x"2e6c855c52924d0bf6909adf5f55bf807ba45c6610136d6ca226b747742af649",
      x"54d3ffd883ef6fd17bb8b257be7536161d8a8d15b32eb6397994d41aabbe8c48",
      x"2c38134fbb1a16cdf8f9b0c09454f9f66cbc9a32fd1c2d1f8e44850f234ea1f2",
      x"50794ece786fb5083851b2cca385961fc20fd429b0c2883bc837e0215ffe6e4f",
      x"889fd409e2fe4cad0d73184a3903f0d2de2e02dc81d559fc8cd9e3b4b4ff72f0",
      x"3a2337477c9a4d64d017d3d56953c467ab53691a3840933730f0130204f26550",
      x"23082485f9fa2a45100b9b330e457ce939f40566657fc4af937a8176f60f9471",
      x"b0bbaeecfe831f1dc005ad9d9ba52cae378a43a61ebed5393e0215175d2fcd48",
      x"b521fe7f11405a656044ab316467b2fa04c660d72419013def84de7e58aaadd7",
      x"803bc6cf273ce8461bb08cb3e528c6618451b73547b026792c93bcbe8d6ef5b4",
      x"4294a49a8b966e1c25eca3413ffd92444833d4a7d7ae74639ab4ad21305cbd4a",
      x"7fe62a9398c7ea5f8219af7136610bf85ae320842fbb64fd47f0266638508efd",
      x"71f3698c23f15c0ef61410985c5c74ea20f32be34ce15c24e0e7f85a56c39534",
      x"6d26345d913c7324b1f27788cfc227ed1547d0bfd711227fc84ca85039ac2ede"
    ),
    (
      x"c27718434c4f879128652de0109ab8ae8aaa103c225ed7fa6be42a1fa20e8e23",
      x"f3a56fb1e72c6edd78fba9ba41ea10cf0491e8c42193fdf39c86b023d6430c06",
      x"ac7d41a4a103c73b104bdd2cef1625b5ee49259a5b866d4327e8366050f27536",
      x"829f29d168bf2997fede572901fd2d2a9d08a9fa12d5a564884fbd23a50902c0",
      x"9736c22e446b92406b3fe90d26b1ee75e79cd81203581001a9e1cf9f5788ed94",
      x"f05ac30ca027a3c7fe3809073c49dc1522b1c189878e4cfdd2be5e04e7a33527",
      x"ddd81b81e2f4397131d6e3bd74b36cdff6b1ce599d4b32ab64d2fe2d38cfdcf9",
      x"62d710c3fff1b5f2693ae50ddc0e96c7f47c130ce4f66b0528093a4d286b68cc",
      x"9903e23b34286c8c9353b1df9071caaae667efb106e3ae40606f37888a7e6360",
      x"09251cb34f6e037fd0e4f951151f81ddf7d9c25f10759badc4c4f9e7d5319647",
      x"e9ed29166558e8a149286be45cd55abc2272fc6ba0f904f50f7b800e39f05e5c",
      x"9125bb2b95a67ec27817cb6969f2cf0c49e51dd9db228944dc20fe201cfb851b",
      x"9fc7ede956fbf4d76a945e3133808f1e40ee3080384e94885c2442946f051793",
      x"a7c595da2a79901ee3d0a4db28570c6d8cce8839627b09c447a1373fae95f0e0",
      x"c783baf180a8ee0f18d5cb476ccd8176bb8c22d9a7ea333d7cdf72b4c38f4377",
      x"f2a5aa5f68e47ec159d6ae1f610f6fec8d5d16952688669c781ecf4df6bfe29e",
      x"3d020713f5070ccfdac7ce60eafe676697deb7d819631e9847656b91405076f4",
      x"1b11f76e64da67a6622ca14675a0a9e67c83f2492020bc9321c3812f1a5195a5",
      x"b7808b4cd7bbb60d51255b74095b72e2bfa1c63cff986f5ce3ecbfcee80d56fc",
      x"09385cff21589396e40ff0c4895cdc8ec445d4f56e9e4b5a2becebf103720ae8",
      x"0e17732fe0372ed597b15c221e869c0c19c4203e910962f5ecc7017cadb38faf",
      x"8bc9dcbc3dae3050514cf4fe7f1389213770d05536740c5ac29f8ca9647ae2d9",
      x"a6c0ab687a05e831b74313c772c50ef9686206f9b10ed0094795c6de892ba777",
      x"c588c44d67d37eab6bc55d0365ac227b7c7088afe4df42bf25379621369729b8",
      x"7e707ef947d8de5ba1731f35606c71385a17ce5ac6498661e1a7941f46b9bc56",
      x"4bef4830d2543339d02092d45418b70e3f1ea27b56d417635be0bc3bd902685d",
      x"60581dd10cca3f1143caf59aeb874cf532e67c8f5ccb28ebc46e791f7284c65e",
      x"ceda940850243d5233ad80a2d65310eddef050321441fddbdfd8da630a8e5fd0",
      x"8e26636387b47de2e91800b10bc3be283f7e4420186bb8eaf8a930580c9234a7",
      x"b0f6a919db22b17e7030f11405e803bf036ca7fed71c036b3e84ff8e030c0388"
    ),
    (
      x"d5da3e32d9633d64e2c875408b990bf07ba613cb8186fd0fa761138f045d1315",
      x"a31226ab2537996fcc8595d41c914e48358c864948edc2653956d6f7e5edc71b",
      x"8fd7af94d00426700adbede960436dd6849d1e362d27c310d06cc5e9d442a625",
      x"7b6c8fe65cfd07f142293ee0e8a0b399691ff0e6287249fdd5672414cc93802f",
      x"9d22cd0b150149ba32cde5fafce4828a50f28b50ce4ed876f4935eaf2fbcbb60",
      x"9686deeb1f537ee21dbd7cd07a2fb7f6d6cb8f20a6a74ff65a149d25d232c754",
      x"6fc89641bcfbdbdf549929bcfed05c9a6907077712ec7745fde530d26d5b7bfe",
      x"8067e0d8597c92744fcab3648481f73015b16911571bfa44e0e79413a13fb421",
      x"0b5f00a205a3fc3249337eb9f87dab09e5fb671daa8792cd663c64d378876fa9",
      x"3dbc7feac0b88154c820775616d55d34c79ad2ada9cf386d50c7446e36917ba4",
      x"f86b1246a362d0b55e042027ae9a4e913ab7f171f44fa9e6cc9792ad8aaeba81",
      x"79a6e420c68ba8b94cdfe7762734878c08f676a3f66b1916fc4939899a5174ad",
      x"02e03da999ef37b9a0617ddbc8400fe1acc09952ccd2ae251730fbf0b29bba18",
      x"4257e4b71a4e74e876669e1bb5ef740c16a717de9aa22f32fa1d7a36f63982c7",
      x"f0399a6c78c8512e200ad550080530404e1ba58fc7c2e848fc21306ebf5d8eaa",
      x"1310a2d81966a9285ff180e6c4f68b3c3c2c292d59cb72e7fea3f998621147e7",
      x"b59c51703527f495216ebd0294976257d1f93c6ade0ea60941bc00e34faf1b06",
      x"e53a17232ee6f07ac2e81f91145f272face5f126697a5ae93ec1c49a444e8539",
      x"994887090e8e6f66559b6118bf954f4da2076380a97619b091601ced8f57e39d",
      x"5ac81ef574b41be010f6f8ee1c0b24ff1a86055db0115574d5833b97c5b00c9a",
      x"2e3a19d310d51e9c246fbb94281a223684455dd6810881d5c5fe8b7ba20fa8ba",
      x"78db86a0cdd66121885e125f43d91b38b935de4c277c768201a44510a93d607c",
      x"e16923c83811aeb8cb54e3c581958cf77b8fa118df03aabd916a2605aef982b2",
      x"0881b1d80f26d84019a198ec1dd8f89381d3cd9d09f34e38f5298f893ce3c110",
      x"354b232d7963557c088094af696232f67eb3c4ce2dd6df1b55dc778cad48baaa",
      x"d89404b80963214fc45577dfd155fff7667596490302222d0558e7c0fa1ab273",
      x"1b8b62113b498767f001fd820597ad199f59e0d5cce39912b3ac60b54a825160",
      x"931acf8a5d1f047212b8f059d0ce7426bfc7f33846e080a9dd189673b1d828bd",
      x"39ae142894b6fa05b6c6172cc6d537310630412ae46ded69fd562cc06832bde7",
      x"ecebf6dd50a68926f6c7419da5b8c85ac102ff99e52d5889f92220ebbe8bd4f5"
    ),
    (
      x"9fad3d579487790f73b773b84c7369bf9955aabb6e186256bfbfaab88baa9e8f",
      x"84a2e73b29dd0071ea801b87160cc40834af443987c939122c438176c4c29c97",
      x"9eb9bf9b9e037e98b48d0a8b31de63a508d2d1ebce806f2b364204bb27058467",
      x"1d39c42959360a120c67c09dcfe7058770fac581e71752c57f865190ab45938c",
      x"368001737035b3f96cf37897b8c1b1cb5aa0dfd0b5980bd15fbde70335e2fa1f",
      x"fda77ccbc69e4f1d8b1e75a9c3b077fb30cec6a04a2ff149028f9abec2570705",
      x"0fdf332c736572a68ae00e3a4bdac22f5f79450592daef91aaa03ee040ee1557",
      x"0c0631464b75e1d506e3acb03ce095793f5490a257b1f64b3a41f855e870aa07",
      x"02041364a007375b225c98a5c8e89c4eb9084ac10e03cdb42a51967e8a6f9d28",
      x"88f938c0001a3d4e40099b5aa77f2d97ce36228ff1fee981908cc94e75f6c8fb",
      x"76ae3fdbcc6d9787fe90ef1a83e6b40b3435832ce51edca637eac7344fc84234",
      x"51c672766b88f73042f1c3afc76c405c3f28c973894bf08ff72ba9d2fc9db451",
      x"c94d3bef04a0f6f603a6f2eb9aa80191af3763330791784273efb1f85e1f893f",
      x"ff4b1d7eeb761c61d4e141811d53faac07c1b408e1bf902e1564ae6411084410",
      x"aea019d2c9497bb9ea2fb9fd555b7cd9870698f5d6ca013ff6cfe9a45c12b598",
      x"143841fbce333ab91c2fc74a90f02bbf51fdff785f3413c8b0d0c2b40815c83d",
      x"53bbafde46793476e537dd75b2a5e791db4f7caa9beda7f07bdc8a6e31546067",
      x"97d92752edc17a0a84ce0b07940d1fea75d3ba150dae7f3056edec037f4d65a0",
      x"949c64264106c5b9f7c7c49e8b627bfc0567eb159600aa0f6b803a962a7d1135",
      x"41d843b25726b17124752e540fd9a925d7d9184d333b5c950094dad72e4adae9",
      x"6299763bb1460e45cff7fd69bd65eb4ae31b1e28c9cded214fe91b8d4ca1dac8",
      x"d7bd89f15495417e342ed9ead343e6203a3571e5d17ef88f0b89ad0b4d945d48",
      x"db07ebc3fe9cdf3585d2696d7c99f6f8c209cb77358bac468c4c0af0440fc0ab",
      x"de549b41c7ada96edf6a0ce8948a95e45a56b726ec7e7ad2c6957e0a14e744f2",
      x"4cc8de3d4a3ce874826131a247ea4ba1668a076e4333a2379e12ba349dffcd58",
      x"647c97d2b551f0019a7ef48e623c8c060d77778113da22ffc06a2ca1cbf8bd99",
      x"98cd6f57ec87d8176f90cfea203a6655710b5efcb2c0ce79688d6b38b7ff3d4c",
      x"4ea4f87e0aaabbc10f03828ee75d0c7278d9bf8c0c03b627a99a78862684f051",
      x"8ff64104262820e4dee0a086d974b683274ec6f2b598a226a4a41c0c8a4069f0",
      x"5a55f2592e882b3c6cea17506816ad2d62088a85d9a61c70ae392b5f8c0c1f98"
    ),
    (
      x"2665391e672ce88919894686f9629ef150723865fdc3a7978d1c6a1f5c1fc140",
      x"ded66520ad5aaf0160915abf3049ed19459dea90de3f24d01cd544a5be1c3f3f",
      x"0ac0a90c65df3386aa72fb1b811e58a8a0ad1cec679a4b66103d2b607a03c275",
      x"0e643725be8ec4872eab429ae5229c46d8fc64c2e38a4a176521dc1b54e0c03b",
      x"baf8d9ec280b85c0a3c3104171b1c549c53a7457c190388e4142566cbd9428a4",
      x"447b3343ebb5dd69e8c97f8712a7a9351aea5422df7ea2d46bf5d0e2f3a7552f",
      x"43c290725002227d4bc4177fa934868fc80189b39b051376f0b7a925bfcbbe14",
      x"5dc1ccf2b2c632ba1c06baf50dfeb6533dbffa1da6fcbcb1a33502f07f9c8a24",
      x"addb6913ad94367032cde9c813bf9460fe6434c7d7b9732e13b25e065314e0b4",
      x"9a30ceff9e022f8329185d3d419d8a1b501d3fa73b981a42a397dfdf576f8b36",
      x"9edf7913e9fab296f4bb867c6ead4c98821734f8a68c05d49043f4508f891a05",
      x"b54d1f0142f3d71020a8b4bbf4d66730df9952fdae2fc4e28b3d01baa79ac427",
      x"382e5f56a158097f193807c656170d9b89efad2b6bbe71e6b1796fded97ca20e",
      x"18e4e473fe95e8ac8ea1a380f3b09234213c32f4ea78bea2466576eb752ca241",
      x"92937def14b3ba56a261b70114386d7f564143315e0e89a664c9ecd0da98d291",
      x"bf51d6ad3100c2b52b255dec347e2a2b3aa7380fd47d9b114ec08109de74946f",
      x"ea3f68697dfcfb49f1998dd2788d58fb0436ea075b1b43c783474fcb8bbee7a4",
      x"b1976baeb39b3d31cd2c674e366f47831f251de0c1850743058e8f32d97fcd27",
      x"5db4b214ba7a8796cc305e1d6dff82fe0c13ec65401610676236dabd6fe6c3b6",
      x"be571dacd82227fc65381ad73488b66d04af921d72c4163cd1f08dca8f5fb565",
      x"b49a7c49d521534ded3e48836611b554f00549440c74ec6833dfd366850d9f87",
      x"e5109abf19688923073b4664ea795cf06f93c7d2f8122ecd0c88a7e2ea28883d",
      x"ce08ad9723121c54f38b05164e22c69d0ce1f594b49943a9624bf7cb8132a3d7",
      x"0bbb65b3441da2146a2cd203e45d7d8bb7b9ebafae6bb5346a226a5cb1d492dc",
      x"4e9898fe4aacce3bea56d48b9041e15bd89f483ac1b0052cc2eda5e1390fa22a",
      x"48321d29cd8a3b4750f778bcfacfab3695d40e690730e41834ee7dab05e9d494",
      x"b2a17a7ae7ffd9c84ce0ec6014ec41555f657947fa1bd25444cbefd6cca598df",
      x"791480bfa983aa7e58a88ebfb8e88219217d918b6d3431748f63c1564572e158",
      x"559e4653c9b6ddd4d0944b05029a66171b07ca9347a15c49c7d032dd7b0da7d2",
      x"6199c5288478d4fbcc22f5ca74d5cae2cd73f73ec19e533a0f4464b670aa4447"
    ),
    (
      x"273be703a31223440066fb7a9f0f0aab9c2805311cbd974a953d16fb316d83e4",
      x"e7e440dd1773dce42b3cfd2f7057704145b334070fba7558ad7545acf09c6eab",
      x"08dce157cb5a2d6cc48e6a49a8c95d8892cefb9257ff3dab734fa877cb228c3f",
      x"64a3132754a6032c652dcca2a0116164b528dea918bf06dfbe518a7334878d5f",
      x"71bd54dac5447fdbbe5d5ae0a68836a67f17eaa9f6b7f15143131c1ad10c8d59",
      x"e254c7acd7e9671f9257f66c3e1fc2fd098eb85e014729a2039899ab8d128092",
      x"f140edfa8959ceb03ef7f7f334e981ae9510e0fa74de1df2432147ed5565f9c3",
      x"fb094feae09d21af5a1d34bff4a6f2c099332c98bd5ca525136114e90751aa2e",
      x"a7304899329cf668c0ab4bd9b56b24f0269b8f13a35281ee42c14bff34731799",
      x"7bb4fb063261ffe2d340ba9370d6029973e7f50d98026dc4a26742c4210f8501",
      x"bd26ff6b54e5d1ed52d8300e960a9ffa17478c548a54ff8bbff03f2dde57b687",
      x"0d6c152effd09659b9fd30123ccc9a92ba02852268f88a29b4d2be5c9743a51e",
      x"703ccf22c11c24af2b4bee6cc8c88467cee568f9aa5b5c2935392fee6917edc7",
      x"87dce489849b434f47e2e0f904831527aed123d750a5770900aaecf676fdafb2",
      x"38d5e470da8ac9c4615e61dea29803fb83e0e4951d786770ddd54949b55735d3",
      x"56def5aa292a1360802a8499fe1673705362d6495058f329a28b079c9900f24b",
      x"b8f393dfb28099d5b5b958f67e0847d39b7192d4238139cddfcbc4b56fd65cfa",
      x"df52c4256d42a29015ea1f697855d0231e98d9b5b919740f0679c2a928312cd6",
      x"5f75ff71eae05800b1d30785c15fa13af527a71ad3a0dcd94691e6d0b5aac6b9",
      x"335d3409f0161d6ed1f97501f6d24c269760cd61514262779acb87095b4ea62f",
      x"5e1f10b3dbe94eaca137a87364b5a3e382a80388937acecf5ded99c4f25ca756",
      x"6a87061431f84c873dc72548ce4fbb6c5c805609ef60e23fd3d2cd5ad6ed9fa9",
      x"0836cbc2a06f5283350e896293a795511dfdaf19b7480ff7ed2c4705726a1da4",
      x"c4b1b6460c8784b0654104dca1694cd7ea65daf941d37dc8bc539a21b7cdaa82",
      x"74ee22057204295ccebe00eed1e2de0f836dabd0216437e7b644c56658adb17d",
      x"dbd7c0a0f44bd5adfe309bd67e9be41d7c4de57f27d0e95752d36e3f2529aee5",
      x"aeffafb01862eb350fa1bfa8347cca8324c4d6137a1f3e1859c9b5df4698f04e",
      x"bad19ab1b180b63ec4d4b01de442fa979a383441b5857cfcf94fb19c49d57b64",
      x"fcbdcba52e441e200205dc6d61e96dd9b5771ae1ea5273b0d4f604bf10d19721",
      x"144200a7c5dfe265d5a8a87a9369500bb956d4984d1c3db69e5950d795be1187"
    ),
    (
      x"79f3258dfa3408f9b4c5d64625c722f18c1e553c870f438a848b12c8f391b07a",
      x"d967a9dcc177b9ae51eec39e4757679ce588f2300c92e459c83a679744d672dc",
      x"9b37537b2b28ff89cf3ab52a1323a21bffa85d9e7d283ffdeba7f1327aa66190",
      x"924a6799020d9b76158fff3cb81bc9e6e0a94712166f77d09856bd89a4b6f50a",
      x"4b87dc399809df1acbe4354f384149bd8cd5a8b9f0c0191a2eb5471f833f1bc8",
      x"35d9635db7d368bae649bff508b509fcd937a2241381b33ef0fddc5cc742d9b9",
      x"76860ee6081cb8efd1da272a44e6b4554e7b65b09dc1fa2e21aa7e766b727840",
      x"4b4d925048362ed0dcd4016a631d0a109b252e78c6c58f13e7438869fb0007d5",
      x"8f71a0aba5be57676be5fb872a6bdd59b766933d185b67b5933216b0a39d72d6",
      x"e26301b9a923933ce4d30f05b0fb3664a0ab1b14a6f3dfebf6aa77de782fac80",
      x"38ad40b6271058a4e81cebda463c7277eb9f7183c79ff33424829f6d8fca3267",
      x"f6b1cbd6f7168a452a9ae0a81adb675d88d792d10eb54bc0befccb053274b273",
      x"88b5cf45df62ae73394d2c90c1f57bb9f11f989fb435c1cb75f8240c792dbfb9",
      x"993a2a3bb554a3be57c5b0081bebe95dbbfc46c77644973c1c4b6b9e968c0eb6",
      x"53a08a4bd3bdf0289edd8dd435f17a7c2be0bb6161d3f0871348ea7b7f26a9ee",
      x"eaa3abdcb78ba5b754f5a8457050f149d40f6bf551c478c9e8d43fd469b39ef3",
      x"83ba3f4d7a14afab20d7461499bf10c1c6832777727183a759d4ea43b6d57c11",
      x"7eb3c94dcaa129e49fe147cfaafca5e3c51a0946460eecba8ab90a69fbdce42d",
      x"ef262ab61cdc32b466b566a50cc2b671d55d056ea2ed2a4715ca7b8e6407ada3",
      x"9a8dd7ea7388f23add65e0626f04477e7b8a9bd4c5389a68149d7c16e1348c6b",
      x"7f706d7492718ed8c1f081e63702e99744d5541f4889ab19f51fbb66272bd696",
      x"793f990bf3bbaaa95c09f553e7c7bd8e3c18dce35337a1062bcb815483bf9e44",
      x"6cc9e241da948e0da757e970fe58f7e82729e586c1514f70b670b2ce6b402e64",
      x"8650c99b4651765658c6668450e5e4ca56a6e58a6b10e58063d8852d30eb0c71",
      x"2168ca131b6f2c088539292af9d1945da66d9a3daf38ec5e79a2bfc240dac20b",
      x"462e3a6475dd3bd460c36bb38b7e4761eac989df1f3fc85f2768fb46cc2218c8",
      x"054943e8ac094ee8df527bd8bc87cd16a5159332f66771ded50452b8ca9838c0",
      x"a20e2b837dc78b12b53b4332c07d11f67a93d9bffb3cdc44b4c3f84c2a9c00cc",
      x"680a8cdf941b6e9935737014e5893c9e8ead0e9f4bed3ce8138ad22a5309e21c",
      x"9e0d7d23e5d47bbdeb7962741bd66d1131468738aa4558b6d03e7cef8913f8a2"
    ),
    (
      x"b3b3873a8ea8d6591f9eb557d131674e5f9ebd2312f8df59605c1381b0232c5f",
      x"18e6a2ad9cbcfa0abc30462a2a26dba5f6c8ddf34f81c67fb7d41867b0fbc3d0",
      x"3904b9887fcd6456550c2e5e966d3f66d2ae1bc4cbb85444a5630e7939e28d08",
      x"333b52e5ebadf382484823fa65a34c7923e7a2a4faabafc7e471cc53ee86deda",
      x"6733362e3d6013dcf14b3f401cb666317a06f99af7f49a8fdfb99fd0a1b66a7d",
      x"1184c3cda0626b9b19ee71eb268db6ac08bdc8704341f971c92431f176551aaf",
      x"a76bdb0d054980495633a074a4724eadf56cd090a78a09a1973d3b3a11b2cf47",
      x"b0b7c8fac6562a59a1fb49c6584d6eea5d1141a7f6aa96df10d360f82df37d46",
      x"4189c725a97d67df715b111d9ac39ce4d4a234d40c372122bb78a350f1add4ee",
      x"580d6e36abf2bf97be6d4fd8b9e6d3355e63911814f8448a928e14ded2759ab2",
      x"b7b210c6f8b127f437b0b12fc6bf4ac88ec6fc283d7017df82fe4431b5f811d3",
      x"645a2ef598ceb79ae69a5b096cb8e3412408822f3c57e0f1970e359cd520707d",
      x"477360c48caefd568c554d574539b3b866b0c20fbcf4463ebf4b9ffc74675698",
      x"7ba3d74b0e447dd24730512a42de846031fac4b7a412fe076104a02bfc66233c",
      x"9e99b0f255454d6bf7b47cb208e6788abae990ae4194df13c77330a2a720b19c",
      x"4d08704b8b026716773694e0be42a225c3ec650183ae351c8bf3ddbd8ec02120",
      x"5498f7534383ebed25eaf6c31a7d4e88e6aa32f7e938d759bb53e2084def2316",
      x"132cd43545d7c5d72f9f0456e94b28019fc32b2894329b7a75923df74d8462e0",
      x"8b00c77aa01fffd94ac5f132784d1504d6869dab4268896f826b434909098519",
      x"b13adc51d9d2b58f876b43445b1fc72b83be18d8f4702828ce64817f3c249862",
      x"dfe23ab641e777b8d2848c14a02c49155ef2fce4cd164543135650ff541a0f88",
      x"eca5a43c205b0871c3a4c9c7dab14314f9d5c35eb8d4aa2833a974a7e6313c0d",
      x"9c9fac7451721b66e38c54fe28c6e082ad06130765b610718cd0e5d8db456c17",
      x"13400b4077fb61357c0c5d4e186f677cadd0decf73b13c919118bcb056f345cc",
      x"2f8dbe46df41d63b86214cc352d24c8e44648edb5bae8a56079987609f9e005d",
      x"c474a183494b34faa69dbf39017b12b3e81bffd562670b538dd4b871b2732c98",
      x"5a98e8b4518588d606ea3f47390568de216370e427885e10ee974daa2ec82021",
      x"d5aefba35a054132fa506ee731a24dca0e6661e55b86b10e1363576683f36eaa",
      x"8526537e3933d66f6ab25033580dac9940f3069be090615af461590aeb90086b",
      x"6b71fd6dd8b2ea9c6d447d37193cbbb578f7587cea13ed36e4a12f89ac22a1d8"
    ),
    (
      x"0f280389a381ca0753eec0ce0b6c3ab4078f12ffbdc57230c577acdbef9441b3",
      x"0bc29bb0fdaf4a012c06280e5306ed69962c6ab0a57592d12944b8466b9a4c83",
      x"5923062e45173aff001567b10cb1a1680e80c2ddeac7ffedc1648819e3636bda",
      x"ec19b80e0a4e09e90ef1b8b56d8fe1634844a1bb7ad27c6c6e71bcdb5c84f0a7",
      x"723442686ba2335a528c29083328d374ac6f8fb84933879bcb1f7db63eae9d75",
      x"f6bbe331625c85e881b444acdace6efdaa5b923e2ad6b5391f533ad0395deb45",
      x"98d837a11ff99edefa030dba4d7baeb7929dd9e24ae6ff7f90b4440882f6deba",
      x"b2b2af255bc82f75305c729c20f85238c0a7db890d0f7f634d6c489a36c14b5a",
      x"d44e8fba934dc433d7be6849eeda29d437be5cab62c4cf0ab1a7e4aa7d3e782e",
      x"46515b895f97360421347f526a68eccb4c926c0067b2fb5a1ee5b33d944b798e",
      x"b35a068fdc6da09e3cf8e870b606fddd7d786e102f354887f9818a1c4d45d736",
      x"1434b9f8f6dde03163014a80a61515f877402fc53c0dc54b4a1ba267092550bd",
      x"cdaff56693d85c81457d0a5f091b1f223c06306c0974af130db7e5dbc21f5a6c",
      x"a3c175d0cd5a2fc2cf40cb63c1192a9c9c3c4c8e8b2adede39f70f89c6b765ca",
      x"7cecb817382f92a2f15f1fc1762e95e23c088c082782927971f76f0f71baf8b9",
      x"0d74d4609d33980a3846620aad918ba17b33d5626753ed48014b576ad84fbfb2",
      x"76c2856dda2dd6e04a56afa0b9e97a9f351c86fe04e44d131a6293686217d7d0",
      x"daf5bd6eee8367071ce4272d765fb864b8d7ed6ae4011fd64d13e1779337ffc5",
      x"56e9f2359b185a447c7c82288997ede1133fe612f953e9b7b5e3cadb020a2cbd",
      x"45e3896b36c173f74a6200f7d36f0c76b83bb1bf9d9b91ea6a91180666455a07",
      x"70e13219ea3f772745e80a7d660e667c293914e1d587b57f1098c8c6eabb56ef",
      x"48957c5373b98503191e3cdf0dd7a0d58a54a38afbc7a3160937b0c0d302ce03",
      x"fdc2200e33657701a649e4d5230084fee4ebcb8cc029d5a68cf43f81329ad4ff",
      x"40d19064b8ddad9ac391a0b3d4c87b897f96b38eb38edacedfc327baa1f9f92a",
      x"05a2dccba738d797d7b4a98cc323b43b5c11dbc332f1942af0ff4495385b1fd0",
      x"4d9db905cb714a914aa37197481f8f4386c7474cf366bc8290ae04f498ebdcf2",
      x"dac0d1b56d498d472c37beff747e001a83a2e96928018adb33fc8bf7853e8d4c",
      x"f8c1c28cfd235edc7e7609e23e21e9fbd79841bafb4f1c6f1a78d62eb99e7a7d",
      x"8786eda5b91d6701e83d4428d0848d7263e026576c466ecaed02a2ac04e651cd",
      x"5797864636aef76b6c2338761238c5e443a29e454fa92e4dcdba4645eeb5ebbb"
    ),
    (
      x"98036eef969c7d99c2fc73b9469d5b8f1152aad1056c5349657c16b105f2eafa",
      x"1b383bbb1de30c91c30ba0d39b0195ed9403b81223389a9d5a2193e84b61b2f1",
      x"d20c9be3272aa65a35c6c4105a97f30c8e181920724e5cb19ec948030c2c2bf0",
      x"f86b359d457837c9eb7611d223dc9b628ee15d3fdb46ad4ea1896f5cd1a826e9",
      x"8bc57ae4bce0c776ea71e9f4e0a68986bf61e190ef296f25a5f95535e7aaeab4",
      x"20ca27b6befa94c81299f7d36d884105901db457c7407f074babc1340970a7de",
      x"f66a5d7d759fc8eaf7708a4fac93132739992cfd208f1bb95af527d4c74cb87a",
      x"ed3baf6ef1998cc69ff780a622ee507804895f51cd6222aa55eee62d61a72892",
      x"97b1f0cf6f9b20fe0ba5aa13589ea45f05114ab164de1b769c162c05f40b6698",
      x"9fcf3888fbcedeaa7f24112b7a357bae238805a2eb5fa5490d03b884e0b9e490",
      x"4cc55af56a7d298b314416be3ea63b133456043c427071441dd60b61bee929d0",
      x"eda29121ebd0b8844a31b6bf7146297876d35dd5f5a14c0cf3f059df7cabeff6",
      x"c1710650f57020c73d6236872fe722405e85d8a1e8c7be66fd85f2bcb54d408a",
      x"2397019d41298bac564a953cc622994a2e4831298b41de0669f5a8d0396b4ea3",
      x"ca2a2f0af65639bc15778bbb7c257fc814b8727136735be7e18b81cd5dc461e7",
      x"fa745a1e1d8e1f7ae3487921df9576ba58b7f82dd3a6d0d6a3f6cf3b16ec68f2",
      x"7b54e196ec08c58c6575d123ec28ef685c0ef4462eee979800e1aae154c6f6a1",
      x"3344a8c2b29eadd28711b887a024bb2d9922a284c1eeaf86824bc8749e401001",
      x"f0d0f9a35d1bb3ae63f9b9f1e19e18f9b82f22adaf8d1ec7697eb047883838fe",
      x"3fb8f6c2e065a8847b3f77a42b7428c7b20dfed71d95733bfd4c71219280b720",
      x"f11f719c6afc437d6287cdec1037eb5e409e777aaf51b5e8ebd1d7e7542de406",
      x"d567b9b5db955af1acb5913910ab25ae78c259b86d11174835a854230eee0cb5",
      x"139bc7cff4fa5773c4db495dac1de8e43854897cab4e78bbe14298cf48638c43",
      x"de3529322498fb96d73cfcfb0195698764222311d0f1ee5ce5faffd4b13c1c1b",
      x"b09b3753db009924c73366a0fef9322099b87ecc93c6b25dd4f01129f25809c9",
      x"6622e0ba3274a9105d462f9034046492737b833d2992f64aa5381eb8b443d4d2",
      x"7bcbeed79880f44b38edf68be621b22d8e17713ed5fafc906ab9b33828f9fc79",
      x"7f7815ec89273cc8e0b99e01d082ae45f34c170ac28e85a3903106b7c021e154",
      x"9039908d890aad5b89f030138ac5c92e584835af277e3cb4ebf4f63b257e3d6f",
      x"90d0041f934966fd760eaa274af84a7cfab03176301748e786e245454460e4e9"
    ),
    (
      x"b156a80739a5dbec08818739b122fda03c4c34088ef0848544b8a591b44b4080",
      x"044a045de1a3a504acd40f09659ba8ce57f2bbc940d69521e64d61fe4ef73efa",
      x"3819b5e4cf1fa7a83d84141c506cdfbee6f20c8a8e619d3e3f74c6f4da634ec1",
      x"f622eefbb08232e8f9f0f0d6f502520ac1fb6280d1d94b335703833c0b71230e",
      x"c5c75ea7c748b9aa964560523b4eda5cdd095e00a4c95b99884c813e9701f741",
      x"b7e690739d76641b55b724c5819f94cf7de21c1ce9c4f09a6d50e803509085c5",
      x"fc0ac3cac393114d68e830c8bf9284864eb8035da518c5c4403cc8683f0236e5",
      x"cb7cf306c4c2b7876df8c2f64c6ce48f3fe58b56b6f45350a9c366fe7bf5edee",
      x"cc76887d601c3d40a44f37305912d2ab48c4af97d691bb9476cf7a336fc25a9c",
      x"2afb4a809225da24e8bdbbddb73804af443b1cf335c9c8f1560a08e20c62a881",
      x"cbab2ede12a424b3fc6e92f287579cf904570fa92464a8f73c22f766b382b4fb",
      x"9350571161cd8734561616b00dea264c9f6a3e9053ffcda4e5337ecc27055d4d",
      x"7ff04c5be327bbf9e9e67d83d10f0a1052ef1e0e8e9e9da951ecdb6b4492af3d",
      x"13d6f4922e138142f5dd38644c6d46abac1a81d333a1b9c782c30e0e2ae75e3c",
      x"304b8f2c1b1c4e56ac74e5832523345b402d3a2f8715ee79104e25a6e1fffad6",
      x"d3dc89854f4a15de2cf525d720feb40455222515d59e3e1ecd5d67c94978adb7",
      x"426dc7e3c70fce5068d48a4227e64a65eead3065d1e99e0b5d572fe48bbf83c0",
      x"368ea85ddf53933c6364186c4d45dd8aada4e8989d522098e6a34c5517edd8a0",
      x"de7ddb7a6b2a40a7e0b47a5a4a8726216d32cedb4e7ed541fcd49e101cfaf29f",
      x"70d46d42b50611f394f3f1c7790cc7e08a832e6fe750ab88ccbf24325b0b5aa2",
      x"7ca78f9781ccbb0bfe99cc4ae23c52329338d82e131d344667e8e5af314e6423",
      x"5ffc34ac72a5f246794ddca4cae166ac58eefa04a3b10ba2f786830a38082cbb",
      x"8746d5e986a4f8e3cbaaed2b163913ede3247c95b32a8cc9d61997146e87d390",
      x"dcd6cac8cccbe1ce2bf8220780f9ee7f130804a76579afc64752d07c96cc606e",
      x"af2429342aa6b0dda693954faf0ef433aeaf18870070be94ea22121e43fbab79",
      x"e9605658499ce0d7e93e6984d2b6dd07ff3a00b746a46aca7b79808dba038d87",
      x"995c1180b87d543a41ceab64ba3d0bd228ba7bdeb88826f125e3f1c9449b82d9",
      x"1fcf950d29c55114c8a9e8140a61d3cbd9eddd2f39af1bcfc8b93a3409660bb8",
      x"d9198cee5a69f5ed0992e6736e32f8714df37c0a6946d0d2fa798508f629fb97",
      x"e9018370ba3689f81a6277ab62aef142805d664d7116d3be9e23738eda071e00"
    ),
    (
      x"e1138eb2ea966f5e6b70e23366f188b38eadbaa60167645d90b91f466401bce3",
      x"40503e99d15f38f804cd865adcdae636775774c5d8e3312e72f0958b18c5ba40",
      x"f639b94f8ea287d7219311114d420f9dc28927a2341421dec221808fe0385aa1",
      x"b59d45fc8295911e08f2b342e6db70f21e9fa5978f303dce69ac2bbd1c0935ec",
      x"cfb9a9b9060823e0805157b3e583ddf3cad25db8b9446b43eb92bb816a52c400",
      x"98ae99c6eee1928d0dca6116d830877b201f214b47847d21c0d1642a33de4df0",
      x"d653aafdb5122e4681b2173fa33397411df9ce7e494dfc2b93f70a47072dcbe0",
      x"5ca513830a22b4df793ccd25b2e2c49b04518c3bbe83216fbbc09d0bb13d8bd9",
      x"726875354d6ef18907a1bbb8302edd634d586d60a726455790e47149659d23a0",
      x"2a87bdd67e3103009e627e3ce5abd145a4c78e173b90463c81cae5c49edbdb36",
      x"23018fb10447731ce30bde97116e3d36a4a8925a882584d9558a97d1cc2d6b37",
      x"d55d0579dd422fed32286d9ffa850487330a30f41a435a1a9d68bfa741743fdd",
      x"916cec394440c92eed4aaf318a9df4812b479059d0d8b57f007323e26ea16def",
      x"a7ac16bf982904c75ea36200ac919577fe8b5b2b5cc89590396ee94763ff74cc",
      x"72688914520fc92a7699cb9f35c115ef882812d4fc66bf2827e2182b8ed19b8c",
      x"28d5a524bb9ded89273a56348b532904fc0708f5d885c984a1d79bdc8cba6e6c",
      x"be821ab3db8701632533f87518a0dec8be988c5bc7476fece8909bcdaeea3c34",
      x"4cb132f3849b03e5474f6ad5d1dc936354d78fbb4fcbfa35d1338ec7d854acff",
      x"3a8bfedc9e67a5f65916a895cf5ca6973526cdf53aed19cd21d0ffdf3bd8d562",
      x"d2b9479d8f31d66ca63ca60c9f9eafdaac304f620e5be919c75c1854690f6943",
      x"87b12cf10d6f8d18cd8b656bff3967c6d11e68d1b1092e074bb26b8c1467f0a0",
      x"881648091e5a083194866ec24a8520aac71bfbffc94e5f2f90d54d3e705d0845",
      x"10410f35644d760abc28c890456de0688ab4dd374c41fbef4e729c0f6091dd8d",
      x"5696eb28647b95ed249455be27572d3e722f94877957259c75681b64ab8f05bc",
      x"14b9cbd2016ad616978cdc3286424412de0c17f4caa0fa72d0de15d84ce2b10d",
      x"9e42b84541d7403ab1d856fa2cf8dfd822387a2220da88d9ba8ccbbb0a03fd51",
      x"996f2daabb3c6efbcb3f5694d5d7b1cd2aaa31c24381b504419f1ebd484c90be",
      x"a765ece560def5c0318e3251fdf296d7881777c75c844079223b19b5912b996c",
      x"4ebcb6cd98a1a47d2a3e3c9d7c7abdcd861bff7f8b4c74d744589f0eb42439e5",
      x"3bea70a22cfc693698ef49ea39ab285caf6870c755d5cb79d93b11e1adc8ceaf"
    ),
    (
      x"411b173d4a8851e049f4b7030f12be5eeb607e44037737ce3d3452d228c7cd92",
      x"eb13fb980d99435c2b11fde6b723a98f8f208bd84714e723b3024d33050c2b72",
      x"6eaf916abdfd90514805fffe0b23b82712b902c5cc935feeb085923def23a537",
      x"c4cc685056b132b9f267d37739713329d22466f106e889062d7ee286135162b7",
      x"93ae6b79ba5218b313801942fb9173aa63b277198b3a180fbba4dce7eda465d5",
      x"3543ed787a30056c9b933b99f3b18a912838b78a474c65b9e13c3917ff6d54d1",
      x"366bb6d42de73674fed0c228c2cfed9c40f10cb24efe7e25bbaba2a3910017f9",
      x"75e8e4503b278698040262c87ca68623e1dbc267301437dff59948e98f5b61b0",
      x"d44c46838e1606d4968756ba7bfa5bb3ff8842f3b55024a401bb4cdaa7e779cb",
      x"c08f888423ff9a6ab0ab19b869a3c579f30db220b84125e506d88412a1cf8ca3",
      x"a662476019ccdb31629971112c772c633d72a776ebbd67db9c77d466f3551e67",
      x"f3612c52b620c2a639f2fc119e82d87b8916ed2a9958cf932a87705c616360e9",
      x"1a45eff2f7555d61750b38e473f4edd4e852915573a136ab4f0b740d2c1047cc",
      x"f2bf566002a3d6375b4e674369ea2825a9b82ad7ebfd79e3f7bfe9845e0d99ad",
      x"7abac39df41637ee0552cae72a12c5ecaa07e66fd9542b9683e8246472f6b0dd",
      x"ceb5f1ffd94bf170694c15b17d66e3a0558d645a530bc23f07a2ee6a7ad518aa",
      x"b8d77d4da32deeaf29a070dd6334f28d17454f59fce8f9866fd1c172f828cfc2",
      x"55b1e1d4bd86072d89edaa4c7b2cf8fd17ae6d23ebb7e968f6695ce072aea804",
      x"7f00aa2539ab7992707f079b8f463aad9e6fcd42708f10bdf54af2584d6464d1",
      x"7d4e88846de23434439f30ccfc00d3cfb749e7ac854d13f7a93624e4e2228751",
      x"57cea68fa231799f91215d4ce74afa9d40ec2bbc30ca433f501443b37e042473",
      x"3ce0d306d916f87dbb650383a11061cc20745c106b252123e8109936fa6b3f48",
      x"1bc8134571fb86aac8162d69cdbaf00ee923cc27b74452979a5933d9f2c8759d",
      x"5df09c459e399cd5d673609f9e3cda8c0838f3aa9eb82706ed623eb641335ffc",
      x"8c2282a25fb4c052da7c96b5adf44f1252d6fe2ef1decaa3b08549d506f467a5",
      x"4b55a9dda60ea6bbda78a2a102746e235d61e24b047637bf89fbde58f2064a2b",
      x"7709c43d79acec92da40595c1840c32d1554d93b3d94c96340896031feef3c53",
      x"4ccb94b1fda6ee9e0c68b1aa70787a5a703e3845277d466918c4444f83b4e576",
      x"d0a15caee96f5086cc7efc11df475f0045c3cd72335f63379849a1b94868b927",
      x"0476a715603de1b4620726b6f5ad2a84c6523158e9f9fb0f2781de9af0ac2a81"
    ),
    (
      x"9867c0c98620e604bfa5d3a9f4929890c8d62b49289000f64f92297688e1c371",
      x"87e1ef22e1c1c3255608f081f1dda28c2bcad8c331010bcc08b81961167ad999",
      x"9802c5e924fa5d81752eec9149e3ef65292983494938ca6dca041fcfe5ada6f9",
      x"c53c02add310756b1c749540e8b30b651d492c4ade45f7d5c851b7d7de75907b",
      x"863ff97904af9018e0e1516a098b3808d7dc072282d3a57dff1bce6d769ea851",
      x"d98d5b645f3171d91aec4fd34c528de03ba151e3057a3b1252d0cefd5dc3ed92",
      x"937dde27b21b6b560cceb30e371e4835d00bbede8443cefda4308743e6166db9",
      x"295b3d370711b4bc1bc11af86dc1f154b7d8ce6ae1743d622771f3f7f53ac41e",
      x"f88937eae892ba8e8c31e61dbd2fc2570f9cd13051a5f3794932dc9eef9fdb76",
      x"1d4055e0b3e49de384d0dd7be714c839c6cc7812d152ada8bdaff7e45d7a9da2",
      x"72e2bad07412c1daf5c79a5dcd72be1b82a5d1725684342d503c829485958f38",
      x"ae7de21343917a884399c30d0a82e8654aa2e524f250b6d56db49d9eb76efd23",
      x"55fe29838b437dce0602cedbb243d40ffaad95e9475835f3b7e5ae83e2e0d307",
      x"b21c22b2a782d32ae2c7835b8fd068b2b497671de028ea0bee03f58bbf637d26",
      x"5272e1d8da40ea871f8cf9d37298c3b48a9e1b61d9b97081bc9fa33a4cbac554",
      x"bb9de74faf2f4b059905764cb9137689f97498022e726c5cf37cefb8b4b38392",
      x"a064659e05ca08f65a24a9727ad4110ef3a1c421c5d178a6abb7c60234966e6f",
      x"c4c00ca6ea205a0a167164280b7e18c022c2208cd0758f1ad94b56d23b30bf0d",
      x"4326ae9541374b2c1de741e633bf7a3ad5dc8de2bd86d1a96d30218484d36129",
      x"0518a65424a509c83821671e8b85b237da9a2cd133e9f881f60693689aed8085",
      x"cc9af007fff85426234e4c6b620b31ea133fd7370db2f98f117f7c5ebf7139c1",
      x"ae6a3ba0225ba7bde9e6f5d241d207149820feefbf84e560fdbffb63d1ae8a5d",
      x"598e3e2115be877e652eb69076a3f6a1204c4b25f30421c118827f696e4851ed",
      x"c355574197c78ea1b10acbd7bbaedab45ddd4b5e8515567aa6690c95fb466103",
      x"8b1d30d750b57437758956e13ca000cbc80c2c66f0e2685f06e69c546d15e13a",
      x"0595bfdc15973e2774257be154396f2e358a3648e33636af28e43ce3c16aa2eb",
      x"0f4d5ff6383867eac4c55b080fc52e21cbf86acd7eea52691512ad5fcfadd5d7",
      x"eff9d9f2ee780ee6bf001792a95e36c56b1ddec9a50c78caa650730ae1fb75a9",
      x"968f0cc67c27fa4e74f766d591f4eafd02d8ed647eb4386c157a10863e11a174",
      x"0e6d77b450cf4ccd98bf42ea374c464ae25d7eb1674efd77a8d325e89bb3b478"
    ),
    (
      x"549ef93e607b2f99f35865a3d02d1725a53f458d78f7c364b105af961f117ccb",
      x"d136bdf4d10333dc42d4a1f443352dba4dc7eeb090dc13b719cd439519a2accc",
      x"2f1e6befc473e5a56c4982c9311748f6ffdeeaa4f177763d7087c2269a289795",
      x"b034a326bf51fccaf546211e6044c9eb9c2827611342deb96783d7aba7869cb6",
      x"b37ce167090ae40cfb5dab6b2e82fa8637412d38c524afc7fa985e3d826987ec",
      x"9ddfe7c57e9a32160d8033aab28c5c84e0b57a6c121f24a37fe84c5c6ca09c0c",
      x"4df4bb8c5281d3232f61a83052080cda37aedcb557f3533caa91cdb4d92fe483",
      x"dd7ba70653ecc48a3a860c28d83d22d1647e28de337195f887557e55e4bc3adb",
      x"232c77125fb9c56ead85b3125f7255585e9e0744dc492169764c664f349aaf39",
      x"e28accd268b5c25b55b25aee60562df675081594b9a1966e6f899fd1cf13660d",
      x"e219c6283156cef432e29cfae5ddb0b285dd0cb905737e7a2ea5a6d664018f45",
      x"ed27122811e97e72fa864d22488d25779053326bdbbcc5cfdaa631bbcdb87dc9",
      x"0f35df7ce62184ca186ad3f93c04659574ec622c6716884c479d462d5fbc3064",
      x"bdf6a16ae19ece6d25c0af41c5bbc21a738196d79371884ab2aae97de9210b58",
      x"aea12964a77227b4b3f6c3a1cfbf2716d667a715e598db8c2f645b797a6d5921",
      x"5bdae0ebb915af48283a33be1cdf94975acbc43ce8b588b2ad6170e7fbb7168f",
      x"3167fd289f818179c07f711f5e9bb4029ce23c693bf92db34e282857cabd04e5",
      x"fe86fbcc4588b46c4920c0f7e7477b5492e7b02685d277fc8399370f54feafae",
      x"063e29876c81e3928b187c1493c67ae9a50381b3c639b05a9a693a8266680ce3",
      x"1891bb10f1a429b64d1f8753a60b3b1b0a17dc0370e2fa09e041c71a4fbf289b",
      x"33991510254389596e52fa4dcebfb918d3deccbb9535c2a284d9bc11252e9ed2",
      x"61aa4e9c8f80dfa61efbaa1fef38530c08eb6fc8e315b96c80d93f3b7b8290a0",
      x"784cd1de32d1558a77c28071f3f2ed8a764ee6ad407206f79c51853570bdcc33",
      x"440a711f8f7eca89bbaa45bee40d85888cc4b197eadf772586b6049db2443e0d",
      x"9256c3d015f52f580d1fe140647eb107f8581f21fe5e326538346788dc9ac38f",
      x"164ecf9e3a0b43c4487b404d6b82d200cc6a1a68a4e7400c83ff3b7bccfc3016",
      x"2a89ac28569c5ef44982e9fe7dfeb4957ccffea4d3cde8a0c7c9dd31358232d5",
      x"dbb80794d1a388e78655424928e3a6dc305fa1fcd57b999d151eaa8d5871399c",
      x"015b6a0e6fd637692ceca96b0cc07379ef2836d89eb488b6cdb8755921138a61",
      x"d68ac287541ba5f0573d50fbd9aa59a70dba1dbd002ffd1a197f2cf7af511056"
    ),
    (
      x"4e263a0b8c3fca31195614271971228dfbad793515cf1d9efa9e8ddf8d08902b",
      x"81d2965ac967efce4207419a575209c41ea3bddce6533270bc281ebc31b0eb21",
      x"ee7b6a6ade8618f940b5a47bc3ad4b390ea51f50794ad3b3b2e9888f450dcd34",
      x"55eb4200036b8fac1dc7054361e4343fcea322b1fc7e604f7f48384377bf2a6e",
      x"e3a399bc409a3cf5d2f89d5668b17543e05378cb0904d295c6a27d49b97cb883",
      x"3d8db47bc828276d7a6e51c03236ea2c19762b3f7261333164402b7b515456c0",
      x"7fb4e0986f743dcac38b7abcd5364a6954ad21619c489776db653ab158f2be8c",
      x"8cabd5d97bc407eb06d3a31cce64891bc01cae3a6d9dc34f4ddce5e943c686cf",
      x"591980c33754015484c980f099d5039188d0a1e73c8ea5940d863e2c0353cb3d",
      x"aac62836cb79ba905193b66d5b82c00b910cf90b59f17efe18ffce5545aa76d2",
      x"b8270e4271a4555b8086ed60e642d696089e1cf5a48f2d8c65fa25400027bd7c",
      x"07c61eba1043ebc54d122d115ea1945e4c06b31f2934363fbce44d85ebf30ab2",
      x"a044b06f63123999109379444b22a1b1224a79878df3739b2b99e69945c5c127",
      x"0614091ff2a504ce70fed88d7820fcc5ce2fd61c95204fbcfe6045d2e35cf472",
      x"5e8014f30a789266517d96da414a529798087931e6bdf173f8e455f9c71d97f2",
      x"ba0ae1d11c496bb3a802635daaa831828e7607002b4790bb2536b36bb7e109e4",
      x"d67389f87ed74cc50e901eda4a7e21d7ee1b4f7c7fc0d0c7598e33b58e4519e7",
      x"4b06737ff6004ad8f20ee4daf48cf18b496df08f7426395abd249cf112926123",
      x"7aed971044a13ae511d1075431ce91162399c64faf9a9d994b6c57936f4969e6",
      x"9c6dc1df7a4be12837e4361a5f71ad892ce4c63a9e73d2f32d10ff9dcff52ec1",
      x"52800faaf5435b0ed706e20f8a42ee3bd769060324f2900e0875361aebf30bc9",
      x"3df6b7fe7d12284124f423db7ce4487eba8b69dc42e3b0230345c152bebafb10",
      x"d3ec1a6dcebc16e070df759cc930a34137ed51feaa3735db155bc03b8e4547eb",
      x"65ce1dae730d0183cc323a7f857747b99cd2307af75e0d7df1b0240e2c9d5868",
      x"404edee71bcb558e43b7cdcc927a85d65ccbe8a7702bd029f1974dd29235b5c7",
      x"950b5b0c8e2570136853e60483543b648baf4e3cb87bf1989e2698da5aac0b95",
      x"6b5fb12f948fa93f82430fc5091155a0b52031029eb1e20446e1bc992a145a15",
      x"8623b283c9660dbeab79b1bdd6b571de80101756891d053ccbbd02127a89c121",
      x"c0d9e61d5c84824d41d929f10d998655026d7ded8d87a53913650116fe5bc17a",
      x"aa0cc25fa03a1d0d336ec17eff742927596950d3c969890b51a83dc5c00444c8"
    ),
    (
      x"bd5c366a377e5195fb47400a29e7e29207ef3289e8ad293c80910e7fe8aed325",
      x"1683fba6a27c66f6bb10e8eaed15c4f4eb4850604616974a29b62b80f7fb0421",
      x"1168b3284010f4d2c341a329d147e1720bfdad60a272903a0bbb7f3e3b37b45f",
      x"e54b570e26b42f67c1bf6a02eea3bd0a246bb31c19068bddf436d746e7cf7856",
      x"3ee9f6837fdb66949949b4670a0594126e80eaa7f8b3b70fe3ace8d4ae8d3a23",
      x"2c9f48728dc0d65ebfd8c27a02806505adf3dfa44f197172ee428be26be15c1e",
      x"bbe60442ba6d6a67cd37505efd28ec7136fd37534de1934900c332f729f0e944",
      x"cf139cdf8f88c660741d1c4eb96d3aa8e25fcec1ce0a8f29022401fc04ae6c3c",
      x"9aab8d8af402841872b7f6860ed5f8321c5a459f9a46208b708cd233036f879e",
      x"0bab0a542716ef5e15b107a172c20d9b19fbe65316ca94888ba882492ef28abd",
      x"656b273896450b130cecd61060cd11bc68b641794044075a9e7e5ad6e64bb791",
      x"5fc4c257d8a2841015bc1ad809821efb1f6011922d238d5b64b3e903db3f605d",
      x"bcc5099d31d8b7205b987d49a6870d4f51c4b744ea221328e71334a8ec3841d0",
      x"6157b2cf9814ab408006468c547886f7c83a54ad6d3e25f2dd98261959af587b",
      x"3d796b8d8b8baf8c47e187d03da28cff6af23d908bd6c93ef50e43b074e9c9e8",
      x"cbf8e221ac1d59566507b4c5f115a6316f7c80e845c5bf6a55df9ab9e8472096",
      x"a6689b85ea28cf025d35b7fc78cd12acec21e9fe972969d9b08632c72ef86f2d",
      x"dd880172f2b422db4f0fcf2d031f06f523df18f17d308e11978203d5dca97a89",
      x"d499c37c4ff122a081859fba003b03e938db4f0dafb27171967dc2a2bcb8810c",
      x"453a110c4e4c88b9f416ae5f4c1f2ab46f4690772ea7e270308be6124abfa7ea",
      x"23685639903953cdd0ee1fd8bc570b2289643b25185fe5bb98268c2d5ddb15da",
      x"f79b61989744100ac53259a2a88255249bbab668cf79e4f9ee74df63681507e6",
      x"683763758876f4a23da6c13da6751ce5fa5bb5d37207c033f8af75fd34a8ea91",
      x"2c40128ee9f76426f8af52834c8f5adc141d833bdf513fc3e4e9f440e1656509",
      x"06c378bc9deeb5c9b313364b730a9babe79ddba81cf80db68a1b28c734b12931",
      x"9867d152276f7bfff0bb2b1ef557e2b5796c84c99df4202146fc57cc5c934bae",
      x"c1e674defc15c09833ae848f9ab59a94a29ef3e1b5d44d320dc30caff134e822",
      x"e51b9cc706d8a3d64a36b9644a58944847dfaafc20de1ed578c0b1389032873e",
      x"01c4b288e2d762f551e8815d74dca27d9e0ffd2f0f9ed3be465fdca0f5dd08bb",
      x"ae87aabb8eef08a7f2406beca094ace704730f936885294ec59559458a614376"
    ),
    (
      x"1ad1076f04ee9598f627e33e0b6fbd5ae0e876e837282b97c8c5de20660ca910",
      x"ffec92b956e6c972c575f3b0c2cd664dda6105c143d40d503f6ca98584d528fe",
      x"f5b1b6011fc1fd44cd00d41b3b05633a5128c503c44d39f205da83e50664cf84",
      x"95ef0289bf677c63c0661623a040b75550262749f705c3aa14361410acb80678",
      x"80fa4ab1a0fb3dea8699b77858e3d397960121273ca7389e1ae8ee82e3c8c51e",
      x"756819e2a9448131416a085ae82150a0d6424a5ce20ba74bd3d2c256b531c208",
      x"3e842459b77db57b10ca77dceeb4e9bc0d12266be166d0a34eb7fe3cb6fda6e9",
      x"1d2b2b7a4aafe77cc493834b4f42ffc2fc74b8576e0a74f1d3cbeb7b0bd449b2",
      x"103d5bcec2934c5a513fbd87ebc2967ec7ad0767671ac1e94a4d5bad45378556",
      x"f92f9199aeeeec0ed1917989277f23b0e23744670ba9ddfd3574207384909434",
      x"5f2f80b4fb3822f1d1e04b8650bf32faca2e14f6010899a34068aa1d3c723462",
      x"27bff025868bd5f3c0ca43f31317c05f69b5fb0b00771e083b0684f292d08953",
      x"4d3731c25ff54046a27abbedcce638a1965d054daa3c4ea3d3dbd5f645e38319",
      x"331c3028456722fc18fa97c80c3753c52fb08e0baddb04b16dca6a44cdf65bb9",
      x"ab3c6af78af3f84a2e089c293ceb449c47fdbb2d76969c022f1584c5517dd2e4",
      x"c40b8be6f732314aa01c8d1b17fbe2bf0bd9389c9b48e6986efc6108ca82edb9",
      x"c81c435bd885f4fbe88021619bb214673d67bae0a0c504687183fe210b0bff3d",
      x"6261304bae3730bf7105c586519c5b21bb39f99ebc2ff80cae7bdfc68132e2ca",
      x"8046a8a7e30729482118f1a62c9ccfec2b6568de8d47d4f27f9e55250715ad04",
      x"d71b18bde0165097f243890dc81e88e33ce4f7d0d764a4c58df5c943c78184c5",
      x"e70bd96c1e22bd652107ba39f9f69f06395b8b9b40baf91e6f96bb5bd786de5e",
      x"ca8e7ee4c4ebf2d0d0b065d21626ca5047865eb25bc88a35b8e0ec410c93dfaa",
      x"e9011f7eb426dbc06d2a8115bf3c5a4a76b338e12b6cc7373deb9e987b4095d3",
      x"826ecd1f29a67e5fb7f7a74f97fc4591d892830556c930ece11df0e1971ff2f4",
      x"88d209f3330dfa096e0357c6650a81c099b7432e98daa9e02461d9ad8c6dc915",
      x"14fd183c9bc7e37b186d8a148c858e2042a865599fbb09bd2b025ce4e46a3f42",
      x"bf7f4056340eb5d6ad3260f792bc1e6316c1745e9142fd2f11399567156850d2",
      x"e483fcad27569e9af50f92a0b5d7b425755d11171b3f3cdc78db1d848404673d",
      x"63608740187c1896f50ca4463cf5a2a6cad026fabb0c47cdae271b0faf10b081",
      x"0dd6543755b984b7cee9ea7896ff91b6fb9791ee7c0f90b4cf127c76d9f30e39"
    ),
    (
      x"197626ed705727a10e5c1f01471849402507ce5730a499f6e113ed264204c89e",
      x"28231875dc10f6afdb8314f125b533a2e9f461ae63cc3c4a72ea3d4c91e1bc0f",
      x"e6ec426ef78d1edfc8ba9ecee4b57a22437beb1c047c3bfeb1ffe12685ceb474",
      x"85b72653fdd2ca2f1ff4f005cae23df66ce3255f950be4a79af35d9756e760f6",
      x"65e9cb48b713da3bfc8d8cdb7bc943cbdce473d8e2b54d859be58ac00396ccf3",
      x"5ce02414561c7f15a61773faa62e490c226577056774a7f9b9a9a52757224f31",
      x"098d22fab6b754be8e581d9d20242964224e8ad90febe98b23e387f378d1b4e0",
      x"fb94937dba2470540dbb5839ed838acaeb6015481a1077ded63e9534be8785ef",
      x"480f7d0321e3c29a326beedebe9142602f207f4e140184e57be57cd83a1924ca",
      x"786ef53679396444598a94af3d1c5a976da745bb4985a42c1f5ec5276962d94e",
      x"554136f8824f2b385b5c79300b645b628b66dca117e58b18743e8860f2f27a5b",
      x"a09302c86da4a75a75899cee29aa9592f35125bba28ae8481fae7998be0ab6ce",
      x"0ec471ed7775580e73ef173afac026a49e098c65daf490524128da556e38cc3a",
      x"ab962999a9e342b004a9d5cd375d49b240e72e02ea592432bd392afb15beb652",
      x"e8f69621555cc2bb2c8548304ea9b85b3ef4700f77a0340962f4c5bd2c2b82d7",
      x"f09dc5f8be6ab7f0f96fd2fc58d7c8a31c778dcbbb87cc072113c91b7f221665",
      x"a24922c7f4c1f3834eed3b8f20492e39fd1e8f85e3db09fa38293d6f417632f2",
      x"0a9e3767b7ecdf734e8456a44786c5a481400e5dd7adb6fde88c82f42939bac7",
      x"f8b48309403fbd7b2977f50635a52776b36a581d2db628be93451ca4dbec5530",
      x"0dd243d8edc32eee8f31c86bbcd8bfc3938ae6f453974c0b47522d9731c21048",
      x"e9a1ac9d4272754ed43800d48db00c935697ba8a5081b3373677f736f22ff9f0",
      x"95d20acd240d998e692893a741d1da0785d14e583eb8eca994c33c5af408ffe3",
      x"e7f544f6c6177ff81c18397cfb6ca34a2f6071d888edf7a530ceef55da1f2ce1",
      x"8cf1349bf8c61788ac778551a13b8b6bff9553e2c388468eaf500e5995e979bc",
      x"ee5b397ee78db11c322cff39c4aafd5b23655a502df9148fb15b3c806a6ce411",
      x"4eca9a7f5784bea0f15214f3c84e36ff357f1daaae1debd9f59a7af88c5eaa31",
      x"6f05f90d6b9b928cf465e3c18f00e0db4fc1c1341d55eb826f4508ab1ba3ca34",
      x"5600755a6a27738d578f2729339fd9eba5239e8546e36b3f5d709bf7263c8ef4",
      x"3f653ecceb84b4170019ff00af486fc03f0978305114a9167f24d10ba47c8e5d",
      x"c24a2a347ebac48d038494b4209d93e9a31a08555ddfd6f9ce67313e932a28f7"
    ),
    (
      x"ef3f5c84484944bf12006ee1e78594297e5ac9286e3b1e0b6012fdf2d0f27dfa",
      x"1500c33877163490a87f006e1a3fa830f09d8aa720ad85176f82a01fd2480d6f",
      x"ff1cb9ad7e53f06fe100450dabb570c6bf974f6abbfaef0aa5d1b6b67a86ec21",
      x"7c2d5f91e4e1da50b2aa35eda64b1794b5a7eba125377d5a0362fbfca00aaa06",
      x"447012895333de2d8c12582e42cda3e87ed36be08283b91432e93ef2b569b776",
      x"027224b34f73f8766833c56cb1831b5c8da877ef3b0c7e7c3c40a512a4011546",
      x"51427b4ca253d739bd87e6b1daef29856badda8fb728f15a2846b7bfeec4f237",
      x"48544dde8745899a754798c46eecbe0266d8aa0f81a991d5fdb7b4d3f9800bd5",
      x"ba2dc42f993725c5bc6c9c30f2e1cabc95327dd6cc8643e75a4dfdedac3c417f",
      x"46042562cf227dc28aaf6ef162a98652b67c902c41235b44591793eb08ab8bb1",
      x"1dcaa1161394f7f5297a55754eb94cd35f87b3f5f60b5049ff39d727bec578c0",
      x"d15a8466d19d2916ada90df91fc4595793f9be00b869ba8b5bbc95b12195fe89",
      x"d7b3ca9fe6e48774baf210f2b19813c27ac7c0efdf9dc1013180798ace91c83e",
      x"01ccde44e9de3c269e7c9beb4a9988a88037b477ba3d576adb0140564b512c03",
      x"83e991d1ff4a21179930e29fbf1602a8b3964640ef2fa126db80d194dc8f0cdc",
      x"791f58bee890a9f79e7a581b96e429444c62d8ee99ce59c13ad622895993e036",
      x"a700cc53c30a4dd1e65af17d7fa6608013c25ef4082ddd60fcccffb1712ca712",
      x"6e38110fd6a3834cbbc0aea78a634938dec5223e55c8d7c73ceb61553e2457eb",
      x"dc31a4972e7066db3436c6caf79c176f714a2785b89290f2e860f5d628a6bec9",
      x"806350bffa27cb3d4d909dd9358862ab45aae78d6d45afcbd0cbe69ecac6c529",
      x"0a1e9243093e3dcd8c520c62d9e021a8a5f862f0d910c4c48ab5f42051a87276",
      x"0e35bbdd1c07fe182f0e9c2b09f50c0be0cc628dca1bfc700ec4d8537e2a2e56",
      x"6a95f1a785fef70b8b1eff5040ddd9195c856da6adcb84234671d719492b3588",
      x"5f1ef9c9bd08f5cde531d21239372644fefa575e86220a8edc88441271f69c2b",
      x"1bc949a54184a88aef899d2b094adb8f783e8a4ee1f4b13c8d7f2a0d1fc4d349",
      x"20ed383773a2acb96f47092fbb31968785e478054fdc20bb636b581dbf4b8a52",
      x"9422bd04cc032ea2999c63fc4caee2e473aadb57ae2e87e98c5dce713fa54f9b",
      x"bfef35fcbe4e324f81ea69b12e53db5dc01cc8097aaf74370dc311cdf6281e66",
      x"2180b6754b9a2b5944506b2c3d13a8a98c805461967cfb210c8f4b198077b1fb",
      x"d052715dacb3f9665c08d1429c799fe6c312fdf7b8d7d8329abd72df8f7c2b15"
    ),
    (
      x"a498b2c16eb7330a17c436ecdb292ab73ba3f10eb9c50c7f650bac86ed6165ae",
      x"19b6aeba4eda996f03aa2285cc0c6fc0adec522bb7921c849fb4e75123daf1a1",
      x"6bf1d5fafcdba9f4382f18a12969e0adf7d8987b35a361286eac79550d7c8622",
      x"c2bbc6caff1c19e27237dfdcc983bb84bd712be40c5b2c49f764aa4581aa7d46",
      x"d3ed75d2ffad3f653a8cb54435c2a64a0c3dd3116b447a46d0af5d1ee38f2e50",
      x"826134a4897287e0fe171f050ef989b95e842eddde26994c652c44700b540906",
      x"586ed564ed2190975c53fb772d4210929a316abc67f11639dd12c71c1cd834bf",
      x"6a3878d43885fc8608cb1b56583fb2fab095f8a607220d3f03b3e3f095a4ea7d",
      x"5071b2dc7e1b34dc9923fdc7e5bfa0733d24a33d69d4f907e229899dd78be3c8",
      x"26835c81f680596cf60c41917eb46065f74c65a0490f458794344ff2ff11e8c8",
      x"fa158014eb2703bb88cda4b403f6dd5a1ec388328722078e72d62807b3a750f6",
      x"01fde50a03cf52ec4598dbe833427ed0152b22b429a9e7e8537b80002e61d066",
      x"1e45e68fc9eec167178498f11bd83b1d6135ed497fc2cba124a6c3e033d8f6e5",
      x"629373deb0e4db3058dee13b6ca1da832a93475cdd3f4addeee1756219cf3aba",
      x"787beea9ac8b9ce646e7869fbe0caebed5df07f56c34a58aafbbafa7634d255a",
      x"ef8226ab28f9063c94202620657c8dffd0206358f8945be1530e263eb8c64293",
      x"e6f4709673870a8abbf2972da27926fcf2b48a35799e97fd5563fa51fe385624",
      x"cec6a8ecdace02f9c81429f4bb28acb2c42fb0ce8d1e56c31419748e142061e0",
      x"de7a064d6c66b4e297615528fec57834a1058f6a51f08bc12fce437c28adf035",
      x"c80719016076eb860d3be2627f3c9d12f6ad393ce3cba22f5d3211d2b92afef3",
      x"4af74766af94f546968cf787004fa98c37c89b737ad57325ccb62f9d28df8179",
      x"35aac8745a7f5744583ec3d48a2425469f3295eef9a07e052671fe10117531bf",
      x"d549c94529924046ef6f159cc17647f7847e2ade3ca176b2c11878fbb26600f7",
      x"c72a3ca1c459a3413c8c503c00fdeb4bb60dc3567cc4812e0f5ed880ccab657f",
      x"2869a4221dc3001e3da87247257c8d46d11b9acdf324929a00079898089bf041",
      x"dc0e58b8c8646c19130711d26e361e2ba6e21709da29a57b7820ade5bc80bd5a",
      x"380cad4b0a4f441a4c10eb7ee38f41919ddae505a577767e483454eba3dcedf9",
      x"6fdb3e9580560f4234a51cbd0566eed3179f0a06eedfc651e0bf2ea0106affcb",
      x"966181927981e8dc62a0be7fd2ca9030409ce5b9c064fe6750a6f3a1e9b846f2",
      x"f367dc10de1effeb79d3bdf668f702bd94882415aa2982b0ee8de2c3d9325e43"
    ),
    (
      x"4ee973412ff211c2b5c6e6decc7e04b397ec1e92acdf4b98fe1391414eac77ef",
      x"2d52980aa56549a164100edca4c749ab6565ee3ccc17e63dbe045d3a2f0e3fd6",
      x"bd552c3e23dd817b44c9e7043077e6045ccff4fc2993fc4427dbbd65cdece975",
      x"72c5a881546939ad692a02cec51c21cc9d5a4481929bae8a810197987b336e97",
      x"4bc7098bd65ca130d2c93af9043b4550f956b8d65957a3bf29f4870ace5876fd",
      x"898f6ed1be83df45a7a98d5b619ca0027600c0b366efadbd8737e9457cbd9f7c",
      x"220be7437c1d5f87c7c273df188140938a28ddba22d1985df79e28dca9bbe22f",
      x"ed32f6109b802d838b87500d11745672b9d7844ab29bac8deedbff4a5a193cd7",
      x"52f346b0d5771982994281dbb3c6f55e7c9f2745f5ba52511fa283cc4d6629d8",
      x"fb16e45a5ea499ef7f45f3b64f868f2268b49a40a88b7bf10f4039af4cdd1ac7",
      x"cbcd0fdd331354cbac81c243d5c2366ba63e67f2c45757ec2aac30c7b8959791",
      x"95acec902c96ec466c5f60c8078d89e69d31f2d41009141af09704e29ea5b914",
      x"d3d4b1efffc10817098eaa2ed027fa5d2a61cbea8daaef65a8ca2c37e8130d33",
      x"4da570a4ac2ed6808563daad39d930053944550efc623f43b412805c7c7b2c24",
      x"59f987423098ee46b3e29c20dbe15c93249d1e9163d125d4b3046caaa4d99f0d",
      x"33921648e9f631a22007588f18f0174818add123cc832f341b7c368a0c28660b",
      x"95d377eab40824b3266e8179708d4016c3175d25a5c8cf7411c7c7d0b86ceecf",
      x"fdd12ae8c8ea8f663d279757ddded08a939bf372d854e306bedac781c72625fb",
      x"77af5a77832de30d548eb30a7c93dee3b41aa137b3449eb9e45dea173eca2f9d",
      x"d4a7c74c25f5259d496c20eb32d63be283e09a89f2537b0638fb2c2eafacaa63",
      x"9fef7e042f562d6bfb063630330fdbbda08cc31c6279482380c5cc94df0999af",
      x"48c0b05cff5206ea9f9ef48e2118e66b85b415e917ed9c0e5ebc479226e60a57",
      x"709098b4a18a6509928c88a0f661353d258bf98160231021528a332f0c2f1608",
      x"287b950c20655a2d442a51257ca49ea97bf766b7bb0b691ae598daa4b7ec0bd5",
      x"07e9af2133ed5d5838c43e0f1e99c7373a6e0fb1589796cb958876d080aed884",
      x"b73e079f1995d082b8f58b4597b5d4803fa255df97f812d942949024f44120cf",
      x"0d79ad4a01081863fd96c64727b4e0532d4c0e7bc320d5c76e6d703505eb0fed",
      x"709e0de3f3c17ee8d7d251ee3fef30eb259f44337746fef16a392696dfec5f3f",
      x"ebcd224773d070711aac8506a437120a552b78161bffdc85998ef4d7d39b6a46",
      x"b955d68a80ef79e14dea573678d5df139c4cda897a096c8b7b69640fdb75ae24"
    ),
    (
      x"feea46b72abbf8af9c752c2c1021fcc5cce66c09ed2d1478c422f1d8600e3bc0",
      x"5483261159f55d69b27522c5ae4ec8b420d04408bd93c4229cd9c7647c4a4974",
      x"6f8c6d8f9ba70f81cb1b756a0750ab52e61247d61b5d244e374945a480e0384a",
      x"ca4ce532c1a0787d1733150d03ae14411f41e9ac2d59b6a6a5b64c01c4dd02e1",
      x"5986033a01fc9d5eb0e8fc35408519af94fb46cccc01d7b5eea080603f19a206",
      x"be61a03b0568e536bed7b99d5046ffc2932a680fbb42e7f655795cd4160364aa",
      x"dfc6859208b4a99475ff9e3ad400f19dd309f146a3c9b8ae984ac51f4c6149f7",
      x"e9caa4ac482198c81823f5ecd4a93eaa720d42c08512a5ec4e80148ef6dd7e8d",
      x"11ec37ca125fc8a8d0edc91899f807c58d6ba0cd963ac9e323faa2d4dd1e4edd",
      x"6bffc7d68176706a4e21f7599dc4a2a54c1009656f839683c96566f85dadd5d5",
      x"33efe7be0f15d56aff194d25ecb7f7f5b61698f5b9927b36d75a1a4d72d4fc2b",
      x"8a4935d616005bce4de9fdc49f3a327bffd885b16a4dc97dd26abf0b55914ada",
      x"78bd2133ed54ebb11ba7fb14e00aa72bfc1b27de9c21e7eb76cdbe8d9bb7172e",
      x"5aa370eedbe615b7083455af3a2487944ff5516e86149ab949a3374773654301",
      x"7f1faa672367ad87e173307648d4e88e6474afbd735ec43dcaba23334c590bf2",
      x"70f1b584f6dc23994ab5a62b734563c791963087573b795954db14e8dfd2ec54",
      x"03f785a85e2075dc243ead24ffb017027215247469e5337bbbf127fe85c15d91",
      x"feb79d5a62092e76cbb73475392ffac2605970d09ebbf7b136205ad00781fcf2",
      x"64364a1e7785a8c558a9a59d089eb53c083ac29d3204d94e637fdc690b331bf1",
      x"9b23c7d6da5c92aeded6dfdaa760a66e32f6f2f35218866cb0707d9caf0dba69",
      x"ce2928433ae27f29524405366cf13203c0baeee81c399052b5cdb24ac0476af4",
      x"714876830a76132cbbc35b02535cd510a9aaa222702be4cae81d339c902e97b5",
      x"006d11a01f8aec2ab59f5840a591a55f4a1338b6e4144132959b5ed6880f7275",
      x"e3bbafe858fb4e9c8c4d9d008308a826f778e230ae7fa88c7b70e42a498ee274",
      x"4ec1aaa101336fa4480b7ad1f265b0183ad5e7cffac25686c08cb95b56cd9d0a",
      x"81370687f65ce4a8ff8e87d3b21e1fa705138ca32bbc7ba858da2002d9537654",
      x"b0b2b203d6d5dcf556a3f62665d277fcc1e6c5297aa949d51d4943fcb2e2fc9e",
      x"72ca024db7613cc231eb1e632f04179c745d59e400e0350039d9335f3b541973",
      x"2af99fad6a0f7c34abf90583b432280670dc99bd2d8a9fd2b9c1028048a95902",
      x"11baed4f848e08459b3f5da01d05fd95a3937bfa450d4bfd77d1139a0e57c866"
    ),
    (
      x"89b1bd1f772b7039110af5d14e110a620befe3169d17f391a44f84a78e566733",
      x"2cd9721759cb4dee469c3e9d6a00efc5578a48179ecff075a836a027e9297d15",
      x"25e5bbda612b188ec8649de6340de648338a910be07720841441dcec3731d9d5",
      x"93f97e65d228ed806267723462b735eccfcbd531e3b54585a92fd61d84ead65b",
      x"2d90b34ec6b891fea85bf37cc449db964318c352d114211497ea9cd4b24f7812",
      x"adabcfd3a44239d83081330cda7b8e00f98f530df9f48f10b1d0c576bbb7d770",
      x"255f2e1aa80376047599b75ab2830862590dacd1c84b2985d15dabaa8c658ca8",
      x"a61082c83b7d61f2eb35279e2b4095372c3c74af806a2e5e06c4d61ae1f6c60a",
      x"5ae2b3a472fb5dbb0df332075f85fd680afb7a3d82fb72bf1acbbae949f00ae9",
      x"181d5e9407be03eea95fd05a9d3e2a387271c7f5c1408c34f19d7404caa95df4",
      x"1b9120eac95b4d3f3a11f36b5b63c786b28c3b1d6e0429d7d47a2f0a9c0f6444",
      x"9236a41f85a27a60180eedafebf707df18c004b13cffe0296308d2280fd66ed8",
      x"1389ae10ae3c59d57f9a2e66212b79bd5e7720fdd764d9ed2c1b0cd49061e15e",
      x"ef0839bcf02003ea8a31605aaa924888de5093fbbd8daaf76f306cee9b4c68f4",
      x"c0dab8cc68d3dfe7fb009028138c767ec42a5bcc7f2091c321c6a6cb641f4576",
      x"f700932947ee6fc1d12d9dec22cfbc35f80beca86770f54906133b04534ebacc",
      x"7749a16eee0841244b16871249fdc9ac944f0fab9c1ceb550eaca5fa88d58338",
      x"e7a74566d0dd9282255b15da8e46065ffff821e1441579ccdd9cefe117728e42",
      x"4b08e1d124b28592548a1cca3e8185be00fa80ade4177e018a4117a35fbf73e8",
      x"4318ae117a076e1749af9660271b9ed8eaf4dcd0c6726e61ca83b9089e60dfda",
      x"a2ce183d52e1e1713b9e9f18c3d33d2a00e27626d9d255c3fcc7e9d62c1292fb",
      x"7c968d8b870bbba00e1ebac84dc61ba9a7111419b034e4e3f571a9cc1a3a5a9a",
      x"57533577beaa29df53b2aa95a009f1d0f78cf8a4de1ef7fd25a5be0c929babbe",
      x"99e5bb2c2749db6315dc948961509b29c2dc0f441340a3a9907d4c3383868bae",
      x"ad51c06dc76ba052a382fd85c8318569c6230089848b3a6ba4e333cb60e159c1",
      x"431d111c99444693840477c0416528cca05a7949616a7a2fc675b3ed416628de",
      x"5885b6b688cd68004c613837474a9bf11a4f181d894e5c485fab767ee1c813f1",
      x"4d75e81e1807ee045b2a85c418b61471de03df5f6880e9d71cef9bef1b9cbb3d",
      x"a2ed8e97d59a38f34614982f4206b8c7e1901d71bad559ea471fc41bd6ef7855",
      x"bb68fcff6533aaa3fc4e6c2779c7a3fd9ed8970668add65cb2c0a4d7268a7a26"
    ),
    (
      x"649f799a7619992bb792a576e9be6939a6cf972ee52f4e56a23abb38dd23aaf1",
      x"3da464e5acf90864b3707aa71603d4a507989a3e59c42d4240e85581ee509644",
      x"3980647231c9aa98e1273f49f10218ae216d7bc428b31a1624fb1563c133bbd4",
      x"dc04ab86788eca13088b381382e26e218cdce659401d21e4c40dc3563b4d740f",
      x"656e39ce916811844672cd4777229f4f791563d631d81d143254bc18da10f7d4",
      x"d21c638115d4dd6ef3e6a4a6b6567d6f4c3b041fb3ce5b427fea5c795f54c6b4",
      x"b7eff51d167ae4a2c82bc59323d17245d824abac4f40d4612ed2f04f80469507",
      x"a6fb29ca8281a5cf94f0831cfb6a1691d2900b4b43ea19aee2fec86bf0f57fb9",
      x"fc3e4f994355cd9977550d5738af8e042ceefd96ffd25c27ec0dd5a205e440e0",
      x"c819758edeb0b90883893f7f09cfbed23b47a6b2465d22cc51cab67e083f665b",
      x"246e252d13b009785050ebfc82e93432e43cee01efeda59c51a604c4dbf626c3",
      x"2aa728a5d2732c0a027bae673fe71202d65be141e165965fc8d7ae3760d37e31",
      x"da2065cb487ecf0d081ae05385a0539b69da704b1ec0b9f3a71b802d18a39fea",
      x"5a8ba7fbda57f35ed83407850a2e8c2ab137a6dd6c5f605b18462ca2e5d5c6ab",
      x"e0ffb68cf7a7c6611ed577c631afcdea61f0a4789137c5189c2d25d4b5d64821",
      x"8488cdfe2a9cf7f2a1d188ca44a6d19c597b22e350704617c54da9c02a7a9a8d",
      x"b800184c65d702a2ffcefe3ef6c0739beef2e0843acb4cca59039117e2bc9b7d",
      x"e267dae2b87f127a0b73c69d93301532c9067beaff5a629a302000a63bb4f672",
      x"3c27e4c5a35d013b8b0e390520c3ff8be7f9f765e2156d89bc8284602e5d49a8",
      x"85c95c663fa6b7ceeeb5d01469e3f3577e4874bce366dc95fd73edadd6305c46",
      x"64e7e4124b5774017b6c434faa37b3fd1a8393b384a4465e8da16e17806c1e54",
      x"e84bd4e2211ef2788e50fe65c8b34e69ad755be5a757983cb2d9d8ba7727e7b6",
      x"f15cd98ed61617c5c5ea9ba8f97443541a7222117ef2fab781ab5fd0d585ff52",
      x"243a809b83385172aa5deefc5ddafe799e75a9597dc641b0a5833e71fc511988",
      x"d8acc56227883e9e6c50004f19cb8118d3c6fbebdaadec61d504ce7e531b5d86",
      x"3e9f779f5a3eabfe4f9ec9842a2528154590631bca10bc694f26576dbbbec048",
      x"d0688ce8cbec353c9b29fcbb18521d53f71215e2eacc4ca1901d6a6919d7133d",
      x"ad631276b516dcadaed0f37e02ab76a2b6a44d167bc6efac4a552a66662cadbb",
      x"d636e76711d9b107e74c40ac27e798b687ea61def0e74d77d4050011c08b0e25",
      x"ec2df0cf50d1ca0129d1c2649da339c01e97878c0fd621aefe0e5a3aa58ec5b7"
    ),
    (
      x"8eff67c59827111f514c2e1c27b264c0756a9932f299028c9dac54e698cdddd7",
      x"542ae71ae7495cbafa171b0d8e34e02053d40e8b90cc51eafeb752bc91d67d3c",
      x"7151f9c36a49c91dda14cfdd304d208c8dfa79ed12b9703cb186126c9c88ab71",
      x"5cd002f7645ce2846e2f5c0cf1dada1224ced55eaf9bb5e3ffdf74fa14b9a9e1",
      x"6568fc04e44e0a079f923f69586d690a14870f7611f6a4c4bcfad49cead45186",
      x"5a87d4b122353914a94d51a52ab3ac982409c9793a5f0a380c72a9acd635850d",
      x"f70b0771f4edd5e430365195c0c32c96e4cf38f1e20c465c2e869a95ea1440b1",
      x"eedece9a6cc31fd6ad89640ccb4d32e7c8178e15b845ba8114eee5a7d79a51f9",
      x"fcddf485ce3e6266a44f56da255cb8ea8866abc7ac73fb1ca05274e9b2138a60",
      x"cff8c6d26572a9401270eea1731e8d57cecee0de49a8f441534f4fb5f7650122",
      x"1416ef0769903bd48507189de008aa5bd4568a902441c57ab389c8749e45567c",
      x"46e576dc38e3b51228627d60e6686fd45570fd4724ed05f1e7cf88b703bf66b1",
      x"780d7db52c1d7af9590765a50f85774a569a2b9b9dac03ae9733cc3d6bad50fa",
      x"d45327cf75cd7bbb8304e8f9c10bdc3c16ce1d6e53c70c68392e3a2c680844cb",
      x"c7a7db553578018a62198937f298800b3de6c5d70f5a2a1681670425210a3d4b",
      x"a2ef21ab66410db9582aa5dcf7eda231f2b37c7bed8bf32e9549a7118912da9c",
      x"a7e054d63aac53605824042cacc75d957e5915b30993e146bb24f6fb33a4f8b5",
      x"ff5b9a50c3e53f206729be3881e0c77ce1456e8f3863f78b8b96c10c9f87ac0e",
      x"6c4c6e21f3e62bc79862325d1620703a9d3d163bf0c17a9bfd4e15299ac10cdf",
      x"bfea6e2be3049e78ff8e7067e7482312fca4c6eea67276018244247aca1e7b3b",
      x"48caab2ac626c6230a81165d18e6d261b212e72477807cf8db87888103559982",
      x"249329654dd959fb35a5c07791baf8d84a38d5721dfc1fb798dd580803f6cfc2",
      x"94175bbe87bf9597b023129014f1b9fdfdd228b8f9901e362176a9df7e53b2cb",
      x"8376db0a15c56ac0213867bf5da6fe8070c92f3b2753db28a1493244dc0cc519",
      x"38dd8465389657f884559362c0dca851924b9f513ba962939ac0118a9995f498",
      x"c57518a190785423828ef7cacc5c3cedebd483739a983b9e239f841acde952ee",
      x"373ac1ff526cc559deef357ba6e31152c378e5d4847155384b8791d0211de6b4",
      x"2237d9b37274d756e2e93cabe87510346685d195f2e7f4ccbf6b1fd74df46db4",
      x"2ea08682e8daed01e373b306ab2743d7020419ee2cd0d005d18d6fdbcda133dd",
      x"ac5ee17674bb1b9cb66ec22aa08380fb66908914415b99628a631fc318de3d29"
    ),
    (
      x"d4f9cddd478d9c400aa9294bd8faa569ecba472f9cb4c40e08224ebf38d59beb",
      x"44d571010eef8baccaa1bf0aea3b69b3c54d2aab7553adaf3d111c7db7a6e991",
      x"8bc836ffcb3c00d1abb8359a2b6280050217d704431f3ecdfc5cd1774f789b38",
      x"3eccd39ed85781307a4358d6c9731c420bc1e0003e7f7be50f5e7d81451599f8",
      x"7a2ccd44200e9fe4988fab3baa13abcdc4601727fe6e0c67fe055795a973e542",
      x"03d2e3a2631739ad642932c1b4d0030b7a335d332aa785f5b600dec7013f60ae",
      x"49c38ce15c69e74d38012b6a8d89e13993850b8494f50e4bb0fe4eb13683383e",
      x"d01dfba14952a91d2561d46d288134ca179232490ee40de214aebefaba020cc1",
      x"1f28f8170632bca7c3bc229bed6d3a710c308ebcfe1e9501c4244bdbb8387920",
      x"8f8728692cd959743dac8debb2d4bf66969423b0a7e158c4b85eac85a49d217f",
      x"90818faa2e6dc71750102d5e3de348200b56b8b1cbc70b13346b7a83c7adf089",
      x"5fd9a57dc3893d98006f54d56ead15460ca517970f80c7c99c40194d696f685d",
      x"90f17cd404b2d85d97c64ec9278714f4c0f23392773015a0db3ab56a093792a7",
      x"ee6188b511decc39202312efea369219e8c7e77db6f5f1cab230d2cc744e129d",
      x"20884b2603762069b42dd5a712b0bbd447c7503a00fe736aca5b8c08fe0cce9e",
      x"307279fe1247b41b29b0892248ef2a727a8c2d8bbcc6987d5889c9c5603a3a02",
      x"6a3df7563d16b1c5b1decca39e81f787372283a03e79a770a88aaa3e58ac13f8",
      x"78df75efc66cb75295e10d7252335ada87236ffe403567d83b295ee2d221fb2f",
      x"a94306101d784817d1d97332aaa7150321112aa1cacd40733bd1b837a991388f",
      x"fad732690f9bb7710e70c6b52934eb116862e3b5ee49746a4171bb9941827634",
      x"ca18ca7e49956a5e736eab64ae433f9cd7141f1aa05bb9d07c216a9fcf3e242e",
      x"5ae49c145472c0951728a2cdcd75f449ae2a22ed6bf96b4adde34a8935db6b44",
      x"0047fdb23dc368b2ddd49b92cb85202100ff0f7e5575ebeab9aae494ca7731ec",
      x"42642c5bfee5971e29ffb38cca2ce93a1df880f7601fef34be683d77cce76f13",
      x"f3cdc51c6e45bc93cf6bf0c84aa5b83e57017daa8a22369d8f18d45265694adc",
      x"88625208063c1ed6bfd8edfcf0ce636aaebb75837052e040d71cb21f562af1c4",
      x"53176f118ae427a3a0bad1bec8fbf989cb845ce6eb54f78a4a1dd25b4135d3e9",
      x"b1bd6177088d65d823fd9e2f7245f18a0223a0aa370c4b4a37ac89c55d5e06e6",
      x"cb3c85f59af8eae66c5eb23933a73ffadc12db38a62731e53111a419efb993a7",
      x"035e89c237fc5b432b54fa6ddadd148b13403f461d3da8ab1389830c00d09332"
    ),
    (
      x"6014ee15ecc62201bd6c1cf9531cfb4aab7551d5d265ddc6146d4239b763064f",
      x"490fd2cf1e167ac89f82a08f2a96bd15efaf17a6ba7e13b192cc9e03bba21909",
      x"3e21a91129566c1de3b40ad96b9fb9945e3641a5e79d9e087352670d56360aaa",
      x"2b847c2bc0fded99f53f82d06783936ce16a549ba9a400a577bd23c1b20de24e",
      x"815d75fc80bdf7012f18c15e5abda251969628b054ea99499b06600737ff472e",
      x"db3209037f342c0a2bc1ef75c5468b8f09a7249de1c1b5ec373c9ea27e3a092b",
      x"9ee56dfcc4d510c6691744a2a6b4f2e181994930ef395297b930801fd2ab28d9",
      x"d546e0427a10e2d2455e5610c8c42874a82280b769362e517e7265824a801310",
      x"9070f9c1eec4da75f4c578c7d168f1898743cc241e0ef04b6be98a0ef547a4eb",
      x"9a5053202878e1ceedd9631338481a6711e8bd1268967249bcf26b06040d5443",
      x"c918d6fd0994b4eec033aa9d5a2b86fb00f4347861f3bc2c92457b2dfee0586c",
      x"f4e2110eb95b5032a49580dcf0e005465dbb8684cdd76a14bce41f007d6a5bf7",
      x"99de6916504c9f3a581470b41855a531b29c7a5b4bfee9767f83d91c58c2e1ae",
      x"c28be3e0446c535e74ae1da45ec7ef6a9520f5787ebf49a8d7d7f7fbde058c34",
      x"9ae110c9e8c407094db8088738a6ae47b53b08b05bc276719f56271622c621f7",
      x"9f64ce0b35fa565efa28ec4897dfa65d7c3370262d6ff4422c77f8c8dc5000a7",
      x"956beff3d1c3d07220fe3b6b73a79ed00e4a8bd597be0122b63fa1cd50dd21e3",
      x"74bb1f3fb052767e672934b6d27e5f8c88ddff3ff5d1feb2486d425eee6f82b4",
      x"4a1192bd2269f916beb47ff3dcc701f3e48069be6d0282ea1902ffbce418f089",
      x"0ca529452a86ce4fb9cc82b4b3a9d4e9a23d395f01ffc6e596bcf1b648a339e4",
      x"7f84e0079f9cdfe083e0eb9d920bc1b09ad0ed76a344ea2c63b904ea274d2956",
      x"63567c209e939141b0a3c1e870fcb21eb6f49301ed26daead206bacdcd370f9e",
      x"8412d180a03076dd3b97ecd85f8154d0135be1f956bae98fa7d8896bf6291913",
      x"112757d5f5b1ab08529fb99405d229ca7dcdd093d5a04b0a2bb9f7f99e76bc18",
      x"d064ff6dcaede8b1fda96bba2fe6fe9f1717f9dc413f53b59d45f2428280126f",
      x"c427a83cb8c82b7356a059ff5658a86895d3effa7f8fcb93d916c4e99871f693",
      x"40afd9ad40a5d473145394bc938db405c7904de658655d36d0ef6e9268035584",
      x"1cddc0fe30e9a59a0155279fde6450109056f514ad21751ebc998a43ddac6d49",
      x"5c71f89849b60b8fc2421b93f861d21b225be060a90e7cf14f92836f78077cce",
      x"5e96c08055f417c17559bb404eb1825e25e1c7268f1ddf99452d44b5a5b8d43f"
    ),
    (
      x"1339e02df46f7055370653aacc4591c7a7496d916ab3906b8c818eb1136a4902",
      x"a4377fd9e92fb5df2459ce9a180bc990d3c2fff5c29447eda9cd6fbd1fbef56d",
      x"350736d5f1eb0c6787f894862ea7dc9ce834bb214af509b93f283a1f89e20e44",
      x"526f084a736493fd265815a8b6e2a2d844e7311add6e142ec48604d4ee0f98c8",
      x"5d802a04be976677a8b84d15505e747e71f18339bba4b72da7f34e168644309d",
      x"2b91626d51218f77feb3c5f164bb64c4b87f6c9c40bf2aba2a92cd9233ada541",
      x"ca0a5b7a326f7da742aa87429cc494831169e4c19126d72eaf83eba360dcf0d4",
      x"01bfd3f6aced3206db6f2cc23124e0bf49bc0f8e3e8c35c0277022364782a052",
      x"9923b53699518232967ade5b83eacd7b1fa31157556a8c4e2efed56212015b5b",
      x"8001d5236c2ad7d2b76acc9bbe16b2bb1dbed7268679fe182bc67803a218a73b",
      x"d1bbaa2d396ff13a9959de3dba7b5e4402f18c95790ddb4794514c5199ab144f",
      x"1879c739eb6c16cf7623c552fd0299a9de0e755f16d6b5dc1728c2cf25e0e82f",
      x"e840ec721f7021a50652a0eb44af928fcd63356299c6abd4665ff43c3bac8d90",
      x"eb3b9e969c1de3caf89d4f45918c8662aef8bb8fb8391ca5a877ab589ee4020b",
      x"48822c4e7384e6e6971a3e6c30dde9760e19f3e83bb2191db0ded9b89a934788",
      x"5db905e7daa209dd1936e18c77780628a971379c2c485174977dd67a60de3054",
      x"4a35dacb49bb0ed9dbc4cd1d9c5fe62c3534af85ec0709894e7cbeb056165d52",
      x"94d8e5d222470a9e3f1681ade18d2ffec9264247f6f9ae955704d62ca47e4b76",
      x"eda7735286a489607bb811d2c682a187fe5c6661f218e512cf0e60c7bb768241",
      x"63481776b95709df2c0f334f12e63e2ac1ee357ecfb05c23bd539e8509b0ce6d",
      x"8f506240a07ad4e724c50b5ab9cc421bdb6cb03e16415bc3a497156a4335b9b4",
      x"f864384506d6161831cda6b928d4524905b798fbc9351068de5cc84d0fa98145",
      x"7cd16bfb417590b8fd151df9c9fbd9f89c65679cc97a1a27bf1269ffac041bb9",
      x"1587de0f4f9f491b543a98f2eeda9b94945367c8a6ca419618ab8edb56becf84",
      x"6a738fac9385dcadded0f22c5f27cd8ba19c608c519cae50a11c08a9149d3fa6",
      x"88e4a681ac206d1b360703dea0eb9e45a946bae7d844bd52400f818130e05728",
      x"615e5afe959cc6d114ddbe83051d3a37f285a9033e5f60e0750e1ffcb75854a6",
      x"83d2cb22b0549efa9b499009a2067ee03582c4950ce2b4cdcdef3117aeafad63",
      x"42ee2c13d948fb7d0769dcfc5a57f085b532c7d6f2283ac915fcacd9463033ef",
      x"d4e8ba620143948ea6c51a06a2faab52dc9775d8a78cacf484f4024c3f4cdfe8"
    ),
    (
      x"498a2ec9f42b695686ea9e680889679ee5d80af570499ba8610f12e99e1b521c",
      x"8e3bed05a4c5955dc18e9244033d16cf8584d0c006fd326d40902bb11d91e889",
      x"9b75cd949ced806e8abc48b75a92bd2dea973334d32f7ae301b8fcd6bcc6f223",
      x"006b8e8935fee49548953cbfa52b61841e05ca2001923411fa371dd0441dc73d",
      x"0cdcc53de68b01d310fa688fa604ae6ade5be28604a583d4d8597e10244ace33",
      x"318708392dac9e3edba8791091ad12b609a3a44adfcca3bcebd8fd38625b43f1",
      x"c47296ad7ea2415eaaac7ea83ac3814a32f69076ad8b0e07445e023f2b3c3fbe",
      x"3de7ea043b86b534ab29390131d28fb73c7f0c837ab43e1e9d3941513e9e1eb4",
      x"512e3b470bd1e331fbdfa5a56eaae547206d4fcd557b329e75ee3a66143c7faf",
      x"6397ee4fe889c3d91c91b25b5d192ee2342478868a89eea98034066d7c87c683",
      x"e67d85849efa6c4ebebe0d05fa354b1b117b5ef3a5ad9880579332055bd33ec7",
      x"5c7485cb85983a199358018263ec3e5781baf1f95c113d08109f2933f3e26768",
      x"c45a9d29f17bc314f2356e38d894b92299b6055f429d6c53c198e323e1dca201",
      x"37dccd4ddf1990355534734270cd476bd6ca19d3e2d7e41781e825ee02565e66",
      x"c4f72a45fd545c48e429c88895dd92889d7d57bba29ce3fce2ef0a124a6020b9",
      x"eedd152d8db959b65d81f5cd3952abc239f83abe489226c91641d57109af297e",
      x"dbec477ae4ec9350ed37731584811b9da7aa933a30ee5e8a18df604cf3b180d1",
      x"bab7898b1307cf218d877f963782deeec4fc2d9d52a483f8335f45b5db2dc909",
      x"cdf45087ed00b31b14116b11edab59dd4b30b13299722fefb9fb6dea92c3c7eb",
      x"37c9b278392f0abe9aa9c8c8837ff5a8217c2d79d8d697c4d9dc170c81e7eaf0",
      x"77e3b8abfa90cfe61ac648e8c53bb222d2872dcf507b8efb58a8a7770c7d99ea",
      x"3c9bede8f96a1b2b4f9a46caab2859ebd270c5a816e6dd6312c40016d5cb9ad9",
      x"3ef09df260d7742d737d8de87daa852d14dda2840c0828c838269df7b13593ed",
      x"62a046c4fe6ed58721b379f5c31ac4bbf79253628c32aae4fc5f5f674964276f",
      x"a84ca07f515f802cabecbbfc8cebb1b2b234ed448ba424dcc81d22fa4ddc1e27",
      x"f324ac75d1c251c260da0b81eeea2a1dc9cf11d96a8cec91120caddc96999765",
      x"fa710635b77af156c9cca2bb12822c16b37f616c0bb2b097baca54acf8e982b7",
      x"5f0ea16b84be5dd09b43b447c531812a2bea7e6e4c93d6b4c1741817882e6ddf",
      x"d4f0e82e9e9f52c393a75898905e3544b1e1cd4476fadbaf02d038c105ef8d25",
      x"7df3c9fb9e70c137f103816e5538c319e973a6cf7b0d73fa9252cc27d995457d"
    ),
    (
      x"22c05106ae333c05e21aa2f89e145163dd30de5530b851ba6b36aefc321e64a0",
      x"fc0a6aac34545f1fc203bf893891ceed9e603bd47b2ecfb7bc6570b831f76d5d",
      x"a7658155cbdb877d6e2006bf46e1f1d8ba32137a4ae1d6087bcea07ca4d88314",
      x"833e05b0a915cd0094b880d6944b5be9ca18f6c3d70b391bc263fdd4807f1986",
      x"aba406e4225f45cf0d8b3107cf2a0a227cd26d1efed9456a5e5db6f7a52e6627",
      x"a36ecca344d71e478d6d254cc38f2640beec5a2a8b3d7482dc63bc9efef73aaa",
      x"66022899a3162f377ac78006af98800fb0a88e247450ced136fce6cbcada7e6d",
      x"cf6887da36c1c2457062255e32919f73b32e85fbd3c66ca777692be96f19a97a",
      x"b8e4ae606e8ab326d55b45e157a20f216b59935592d2386d6db02ebf60a3d19a",
      x"72ded81e39dbfb2e352a5716311d6b50561e842c118a8854a093f1dd620c9842",
      x"db2666360695b76fe31cb5c3258e3a307cc38cad584d72995f74dcd79b8539c3",
      x"1651e92093e8b302c82450673e12e89bf87b4d27ca1cb0c7a65c9a84ec11cac1",
      x"3adaa83ad1876ab7ff8d5002f947e2152b82017b0295ece86797192ab6799349",
      x"551120fa151c37c903ef7a467cbcdc5f6339a621ff9e56d1af85f805ecd40a4c",
      x"941a657d7f587043cd7fa99d3eb2c686ff52d0235050dfd6ceb1022e840de8ba",
      x"ed79a65992e1e0c1f75f5837db2e5ce4b0c56dce16c2bb93a80f311c677ac342",
      x"f987b273851e331778236242d0b0ef363d0bec0b75eaf3b2fc41b6ae74c85524",
      x"9ef09ec2d55ec4fac65bec26f1ac0c2bf70200f7aaf5904544f9ade59eb3c432",
      x"fe0b3ad954e163c0a66e3d52622aab252e714f0040ae45e9143fdc7b320b3d90",
      x"6a552c7350605abb028bcaf48c8fa1a5188fe417eeeef390b1520a1a59371dc9",
      x"686a43e7db558b3d62d5e5e6a4304e4db6068f76c0066bf75e3dc74d18eba2c1",
      x"7b966feed587efb41b6b58c86d5fd9f753ea2e176d125c4aa657d22af533f79a",
      x"f4f74f63d1cea75d5636ecec7823f44d532979a8dee33dacb1491c55f728e98a",
      x"8bd6fa8a9b1cb299e3b8136e79ab8a94782608d7b8f8f950fa0e490d6a94b7ee",
      x"87dc03fa4efde8aa4cbcf3f0121e79960d1a634be2462d3505c0bef88299613c",
      x"89207677fca69fd8fe3d3c8dda52d5f19c992c05644fa1fa96d4b076c6a04ff7",
      x"0af1fa9b142ac84105a842897235004b19e117079dc21f21b748ec36729a2b6d",
      x"21501910169b634a53058cbe534ebc8be744a77ae46cf1c2748ccb1a172bccea",
      x"328c2604943604f07fb4a0f1d5366f868bfbc99b1fcdc9f4bb57cbab95d60bf2",
      x"d82d9338a04361bc3d7c943bf266e11c9be3b70fb57e9d6f8083dfa28e4955b0"
    ),
    (
      x"2aa4d8fd425e6f2327025dc47703b167daf177aefa2851ff39158878668d76d9",
      x"e6770be40a0f0a11352556d8b685b5c545701418be670297b923287166e73ddf",
      x"563ee9bb701dee622db88a6f1e18363f539c7cc06ea53d0f5433283e4b962fa1",
      x"0b6e6d35afbb62af818e7d4bb4c426404adc99b7dc86444710659521d1d6f82a",
      x"aa0ef1dafa8d5479a8852fe801e075ddfc9df4f3e12cf5674ae419d2ddba3306",
      x"045ff3ba19cf8d09b862e8b9ce561f7773040879a105cf86f71364b58ab17e23",
      x"8485a82941f176599c64834a646c0fb853596223455e67d07eb631457e919bc6",
      x"dfecf5293dce71c0c8a63d989cfa3f70809c554516bd9a95cddf56f67bd76c82",
      x"ea86f53175a38dc827d4f178043b0bd4db30b4ce6dd2225e9a4c59a8ae90381e",
      x"974aee3299a1d1444260bd125b23f04cda4662faf90482406fec1fd15873a599",
      x"59cb0f08aa8a11a2c0c757c7737bc05bf1279c20731cd109ab7495fd0836e564",
      x"319171ef070a0664f8364d463ff5c0a10ef4d92996ee221ab72cb781e17d0c21",
      x"fb4e2a3011ea7be5e5ed6776f24219da6f0775d5acfd02de7052d1683c8b9a8a",
      x"2c2e8d2e15bb5f4b7031af3abb77b4e177a177da6cbb1d5932016af6dd243b2a",
      x"b34e31e16b00c4801f39d4627f853d2bd2b086c114b4022bcb4a04d8801dcbe4",
      x"4791abab59e7b5327c43ff852a0911cac33504b49832285ed75b50c3519bb825",
      x"c13081758ce9fbe0a11b7b0df3a5259e7347c431b8eb99aebaec63a5077b0a11",
      x"a48489c2c91e09dcfd5a1cff42161da10d0a854ae92e1f4668fb2e0078f36b2e",
      x"950640fd468f6e9985221fefa4f406dce5d4f8d0ca7737d2ea27d39d12625dc9",
      x"779f39437f26f1902fc3d0f2fa57dc2d3a4a73cff653c948637917f65812be25",
      x"5b8b37cbb3c71ab6f11be99f5f270886340ea74e43559065c77cb41502fc5feb",
      x"48c1c63e47de6c072b33d361d4520452076fcd4c52958446700e41d462273e18",
      x"28ec1789fde1497b91322ead92d725e66588e340cd3f2f8138d2f123be4ec20b",
      x"0591d056e638c060c58c9929510266311bc80fd1a73539200296a549aec56896",
      x"abc52fa7150c7e7fa905da5b806ac9f7bec43c8ca30ddd09298dbbff8dc031b5",
      x"0c986146eb6e0cef39a061816b4683e844a85d58da66b77f4301231848826157",
      x"c51aa573ee8cf4e2ef55a3a773f8902b9498b36bd9cbd88d81ca7698ab0ce99b",
      x"72595f95a92b0bbb3c0248048ac61a5aefd8642af6b4de37adcaf09330891cdb",
      x"ef8e39b2da080677877b0f255c5877c87d12719ffe73edcf7b50d2f10a7eca05",
      x"4a2008d667809bead4dde45d5d2a9f5e9fe3a44f117fc7069b3ae22b89bf2598"
    ),
    (
      x"24fda0c178f860d649d9be9ce51b27405fb62fc78721136353508b6c251c84c5",
      x"d6b30aad6595e30b6239ee75a6ee637b2671a2778067e348aff92d4317e2cadb",
      x"d4a93540e67200cf6bf416562f6314e0c877d7fab806aa71a6316fd3621c526d",
      x"869a8735e6b7b7975af455b76690fe09719b44413b1c08892b21c63f85c93ce9",
      x"021ab0e13c8b77f03d9a6b8160ef2f70f65792fe1c4fa0f3027c09baec347f5f",
      x"0ce1081ceeafea61996cbe71742e4af65b949ec9dde2e3f435687ec9a0c6ed77",
      x"cf336a75810da94c3c9bf9b954d22fea6a1e09f1de42c69d72a6cb3f5fc37d37",
      x"8e9bbbb721b70e64b57eacf382e52a16de8f6a21c81f0026eb99b6525804e14b",
      x"1c5286145f986ca68d2ee3563fc5199416dacb45739c4c6c6e390929a3812ff4",
      x"c2a0eeea48863a4a4a899b9a3340ff41aa6304b01a5e49acb9a5d83a4ec4b4a8",
      x"1f55954a51d92c5c55791c62a293d0ca89d2680c1fc251bcaaf5d5ceaeacf602",
      x"04ad9fe76e6cfd123531e8a91ee590812b99a295763136f8f14a77da8d6af4c5",
      x"33822350696af55862f81f59cc86ff9b98ff66d47bc9cecf5a8f35c720f90ebb",
      x"6b8099f3dce8ab0cfbd9fad93d075ba1bbac859753d19323e31c66e162865be2",
      x"1a6edb1efd9b42012f7047f0e9123683d8f268ff2ec42c4cbed736b9ce63b62e",
      x"f69633a5ee943840ef0c0ce15960a26b4170e8fc808ffca8b963adf1d5adf2ea",
      x"6b80ce6e37d37f8457481e81637d652f196e9dab9b3e6b9371ca5a6e4efa0f18",
      x"b22a3509051d3d32f7d03226a74f5c91a7ee91285a2a653abcb6e973a1354870",
      x"e9bb8585d2e2faf4c172a409bcdaf4eb1425a64d3f4afbd5137712f9c48875c7",
      x"7cca73ae3c4660404ae36f0c5fe4b49d6f860f45ddfaa460b87e42caa14bc30d",
      x"b4999ae06f2ab34606bbfbaa99809c1a36c0f5d50135288efac40c3f46957a99",
      x"0b6ac4be1f382df502d7a486de3bb1314245973cf71f6dd9d5e7edb1d0846918",
      x"ab98de55201eace670a669331ca00416c64b05b024e20569b152b0f6e6310af3",
      x"65d56cf9cb43ec6b06ae5da69660ce465f46c138800cbeaf85180e434483110b",
      x"3cf86f314b57e0de6044e3c6b1fb67b3c41e16ab1cd5dd9c94db18c7b34b40a8",
      x"24f17afc4d240ca7b7f87c77efd2590eecf18b0204638d31bf2b68b9752c4d32",
      x"58cec460ac75feadaae0f4892250af68311c75bc24219dbf4e86e69e908b3000",
      x"b62f3c878c849cd3202eb5c43af0ecdaa6f0695152082ff05402e0bda2432cd8",
      x"e87c433aa682f7b3bbaf3fb865096a67cf8b97e21d4f4329568bab1a4eb38523",
      x"1e8f929d6296a285b21ba8c8cdd1c8d991b456317f28e6f3f003128525a0015e"
    ),
    (
      x"7cc37787a4723e13e7a6825f3fae0ced3f6be1842c4df5000875edf8ab99f86f",
      x"64ef95ebe1e21db04bb756aeef166bd535c49f24899596fa6d7eaa4a3e7dbef5",
      x"8f81bfafb32af6af2feba2b7e14d10e20d8dd1b9118050220dd4fc987cdd7c01",
      x"6e10e69e8205e2691121a8ac3d9ff32be57d1e323de664ea4307a77d390ab76b",
      x"39d05a33bf4c46e12fd8983ab8d3b005e14da8472ea83f869902f58be9435b14",
      x"ae7419dd9872f001b3006d9d4440373101c217c2cd0060ae5035ba017909f5a3",
      x"4daf9d454af03f8d26b2e484d5c1db31df5142266a01db7a954506043e60d21d",
      x"a48dd379320172cd740ee3e9c6135da2d99005a41d42175c730ecaf8fb7090af",
      x"3071704d55565b9391190124a88fb195120b64acfbca93fe74a301bb6c8e86f4",
      x"3884728d5c5f3f976af19e2f9af07dadbd1e9b960dd6b391125a51f8828e753c",
      x"d84fc941c2e52412a2b8c1b313875b3d601850a121dfac94e5e2f2a0ef0e23f7",
      x"bad6c0e1a9fae8e49d65107fa91ef6f18c028b9aee8fc34eb6793c4733795597",
      x"99d2d3006d4a1a30681ff933d4de95bccc53125ba774d59f368e7d0fe8608f4f",
      x"182a4e85b002ec1dcd621644b707e51f9b4b4dd751789578c638274fc1dd07a4",
      x"bee657eb2a556c088286bd60999721b59939b459d871f412a43b6b4289ae281c",
      x"bc85d5d348c2f95e5172bdc4b632c0a3dc5a3b4d2df4b6098e3aec6e305bff07",
      x"e336d40c8ae018dd548000eebb98eecb1859626c615421c2149d84dd1a5be236",
      x"231d91ae29961e216f46cc43b3f3b52fd894dd795a206808e40823bbddf201dd",
      x"95c45755257693a0a3d8c0ba576e6a9e7c854cb9a722a22e68d6d97df74e63d5",
      x"cb4e79a43633cd475b12d894e3efe20a032c0de88e6532f59342ea6dec519633",
      x"e36bfae594727aedf33a19068f3a3b10f031fac48414c36c0812ae5272583e7e",
      x"023e4ebdc2218d8b7b6a5be91efc4db9c1b6e2329f0cccafe44c4f0d5fef85e9",
      x"a5c41a4e96aa72e5a6226556fcb377f60c23843af88ff72d3f09866183fedfb2",
      x"30f6943132fea55aee724da0a7678876f9fc5bed8c7821f773eb7e2945194389",
      x"625a642a6ba72f0a54e3f771e0c2348e9b30c93d4845e24269a883750234edd4",
      x"bdc8fbf0c715df3d5a3863aa9d8ae5b45499b5824cbe97238f2269d4fcac08b4",
      x"8fd7bb2f32cd624a5cb457a281790374e9a0ab9f1b92d9db7efd2e8fe9a4a66b",
      x"5f7b9b3c0859f4b71b60ac8aa388db0beaea312504331c77a953414affcd422b",
      x"49448a66befeedad5a0eb18bcec339b44ea66f6070bdcfd2849013255a1641da",
      x"44a694ea1d7929567a0d29d91cc7b8d617c190490ce8b57b589c915a505ad870"
    ),
    (
      x"792db055695b9ea1448a7aca82d44909308d316b746446d171bb031023699465",
      x"f7ba4ed58155870c4a560b26e6238bbaddadb7b86f88e3c07e06517c62cfec78",
      x"071657f854cf3c9a0d65c9a0bfc8b0aed354fd156b0e4600ce81bcb7467c3b64",
      x"920b92f5b7fd6875a32af9d6c03abeb073a26f119cb51a3597d34315b542408d",
      x"41b514d233ccf94f79a35b1582dae4656499419bd02f2f4f2a2339769a5325f1",
      x"fb5c68ee3f1e6270b4c2787a20a6484fda67254383e9444dcdeac931e6d1d568",
      x"fcf40b1c535c3f9a79eb072d66acc3e14f08198021d2128dcdad86257e77073f",
      x"07f12b2efa62fe62f47d85fbea245383fbc44d7ee9e0a76489cc9c29d5241f65",
      x"36b55f87adfdc15622771edc08f91e9052b49ee5a51026c7fc74c19fd249b6f2",
      x"3d47560c0ec037771cbad299ddea3d44ca452e173b5c623f2b1604faa4da2010",
      x"ff2e882b3de110b502974d3bc3f6046e01fc26e848f1841acba31f555c6760ab",
      x"b1bbb790a89df02ab0488154822d743bf51e0324540bfadd01387efac0775bc5",
      x"d9382f0d820afca512523ed4870ebcc0193e7a78569bef3dad1878d9f19e7f52",
      x"1982e7b9fe1740b6d199a12fe33775f1781491bab6e95cea5f6106f5369cd0b9",
      x"b6ff4351c290f85a1185e0787f7a8028e98934baf2a079bfc263e0f3940f2e1d",
      x"abdd7430c49667ed1fc9e5f2c5e4b4bcb0287d6fd4327820f37c15262317b7a3",
      x"d6f996c15b5875a1b43bacbff6660b6150e7d84e1ff6bef47fdb72c855b90690",
      x"2dd11d7d6439f41a3b786e75558cde5a2904b299afa0a9dfd748e95b206abfd1",
      x"f6da37ef61cf290b6d50bd9dc9abd1c52e15f0d38f0a52b6b9b2710353bff961",
      x"47a58d16c8fadfff1d731cea9dca0b0176b89469d1595076ba4f711f4950833f",
      x"c6fcb7f40ccc29563e7e54f5cb5b9b5b15d830309d41b57b03dff7549370ae62",
      x"f188c203e300953623176f85a88c507c4eef28969250ec0c3d22f951fb2149ac",
      x"ee177883964133a7e39dccff2af331cce4e7cea570f6bf94c04624606254d2ac",
      x"890615ff124617089d6fec34a767a155b59331adc0f4cc7b5885dc8354d0f6ff",
      x"72e6f9df3d6d0ca992524cde60e78f2c07e6fdae7a7871cd3c28588565c60808",
      x"6f313b4b3ec0a4c0f5230588588071cc4fb8c67258d515d617d1665885be48bc",
      x"3238880aa661dcf557d591ca5aa631905a14b2689a21aa8363f99940657e49cd",
      x"715d2724723fc39893ccef354696da5af05f736d4ee40fb926b060aa4ea766cd",
      x"2d16b900fb641386a102a5c4f33de42decb3fd9ddc8e1278627c88831690e660",
      x"38bf76b0b0c73c85465410f41e986020fb31ea32b0bfeb4d5184803e7107a4a2"
    ),
    (
      x"bbd12ca1578c52583fdb39218e134051f6e55a940d8c58b5a21665d85288e977",
      x"97b45e178dd2ddeb2a6ee980f15ff405489fea6c1616b3e076c9f342cb5956da",
      x"144349704882ec218b75ae408314720d2578497da38b0a753535e609b0b12e33",
      x"6f6f106586cfa42108999e8d462730379ea72b83a86366916d162ae0877aaa2d",
      x"0b4a9f63e6051ef68cb22c82e4e7be132c62123d24a8c272f1beb633ec9d767a",
      x"c3363a4f3d66dac18fca9535a12fef2afa651211e53b170b99590f521522fc71",
      x"d39d1ec42cd35b6f2a088c184c419c34fd07fc564494e36fa95dc0ea8e95997e",
      x"3a29e91c3b5f78d20ee0472d595a3e68c38ee5909bd6ac5c9b193b9f612fb14a",
      x"3291b68c8d0c1aaf658b826643fc6fc5d755231953a43697d225c31716cc8a5f",
      x"677a1bb2bf68f02f3c5f0d055209041abc90475e2d0f473ed0b648c9b882f5fd",
      x"1df74112320a220f505e66880c3518b6a2edd7988cde854620fc164b4f5e694f",
      x"442400d50ee88ecb7af90a59a1d2c153bd564c03754a472033771d34594fd162",
      x"e4bff68096f0e1fa7595858beb6732ff4ec21e97d826f4822d9d2a86a73f17a7",
      x"2152fe58fb012f7cf1c7b30fdc5b34d00665ede875721edfb0bf026927792127",
      x"b34bae62bca3c02503c52127ae30d853fce78a773040ecdf58a21d71f47933a6",
      x"d8cf8e56aa6baa9095011d06ab2232caef59251f6a93a55d53eee495f17ca474",
      x"2e05521281175e1be990a804f5d3e16c59d2b1171da28ce0691051fd0614d314",
      x"1c127ce7360a02762077c8d3b3c4fcaea73475341c5ce6bdc649b35cd00ae692",
      x"7a6db14a1f7e69da68b9b430e4ff21176c33cf0ef4e67a93f48a3d8f5caf4c23",
      x"95425fe609ea8bd50c882bb7c84c4d7ccebefb3a7caac2eb114df9c10cd00427",
      x"dc82e2d18777d1874d594cc3f0197cbb2562375002d0850f5b10eb047248b581",
      x"c76a997d256cdb8d2ab2fdb4e4afe4a415ab91adeb3b5518d0ff34aa531b73ad",
      x"5877ae28f0bb6802797ce8e1aeed09565f79dbb4500bfc0d2dacb63a1fdaafd0",
      x"3544bc0f773d5e4c4af9f8da835034228362840e44119c84f0dfd42b0bd55527",
      x"daadec46c27816e3623654905701b50fac5376cdb39c1c098e9f31106c461e3d",
      x"052212e4e0d8052a17ec2b1168cc60e4ded10d921fdbd7f60bbcbd397382d0f5",
      x"6ed50ad8d4722b3192078f2a1dcdcecbb86c235c70d7645c99b0c7f2da10116d",
      x"7e0ce356d434bd53cb2084954740b6ccccff72502fe0b8fcb531816ea5bf71ed",
      x"df2b2bf0326433d97a281966bd85be7041875a56b3c4a19b1bde8e0a198672cb",
      x"75604a97bd9da82661f479ca54f527bc00c222aa93a4c74907e3ded4dd6551e0"
    ),
    (
      x"4089767e649325891a1f1b212a11f7ce856dd34930bb858610046b14a66a0232",
      x"077760eb83da99341fa641346c5b1807e614e3e902491f972e97816f6bada765",
      x"95630b0ea49574c353d852d7067659357d0539eb9b5fe062b0ed0c92ac67684d",
      x"d16a5fc264f150c766e7b931a4a03c130d0f74b487221928ee8f953f224b2eb8",
      x"02a2fc5b8968a36cd85ce0aa2663238266c3e87b14b37ed9cd257113db536b3b",
      x"bf8cfa3ef1044ef53407cb69d7bc67ecb47fe6f5d6242411362c4149b1977baa",
      x"190a23980da5b93ef6ccff96733e1f8d3aafbe57e0017d883823e093517c3319",
      x"306a959ae226d16d510710b48e4f88b6104a3a0c566bab990cc5c4ecfaae5ae6",
      x"4f7762baa031b47e05c3d4aec17f0f4bec753cc7f166ef99ec7dea4e5295a843",
      x"9271aa27c1ff1ab08700076f43a95aeba76a0ba282463188c5941a957c1db210",
      x"b4de95f5c4ba9f4426bf5015d190cdd66ef1fbaaa4c9f4ef4ca0e3735507f379",
      x"6f370c322510bb1be5cedc40c9ca2e694c2b614ac2de0e582a94ad9ca7dfda58",
      x"44e8dbfadd5f4a876edd59d3894d11362af92fca87939312be1b73838e25d984",
      x"8c83126e49aa29acadabcd52a0fe1e3850d1484db17977e57ab401b8c44956e9",
      x"7df2b93317213780afb2a95abc755892fd41d5c9d7c8b3b28b9d02bb9aeb699a",
      x"304530eeb7fa8310349acf2d18fb9aad9d637b73d8e8860e3e9dcb7a1ead99e4",
      x"2a8d70f2d4fa9fa9fe27304424a4071f9a24d51ea267f32f5bce206e0e280a8e",
      x"6eabc44e65986913193c7ba591f82dbeadd5d65c3f85c7904378a3b53fb1d546",
      x"87b15d7fe02d107aa7a2aa529b88e66108fcb6fe1f9b9e89b933bec39aa2d61b",
      x"41eb46c01f7f41c8e5e3b4a3af9c1e3172b5595de1485da9697965bda088bf81",
      x"ddb3c15d7d743bc69a8f2027f04ee5f057e0bb1b973a5d278d7e7f4be051397d",
      x"9bff76e1eb2abc9495cee87acdd91e3eb02e6cae615effe0c6e833057254b572",
      x"1bd2e3d193e7508037af6d1219b94eb776b0fa3108ed1a19cb6a80adb2f2a4a3",
      x"4b03c62b72f0461d24975687932aac0efa884863da0bd28f23998215d0cede6f",
      x"5714edc661ea8e60c470eb156cf24863a70f2ce9a44f30f8b66f60f4a10757dd",
      x"015a841bf4bf2a6543fad9575a5821b20ca2590f5b366471952ffe8eee80044c",
      x"1189253c3630ecd97bd763b919321fcd86f6f8c3d27813e7a00480dc0da62b76",
      x"28777cff57f36125fb5af8e54328bd1475e30452a407aa9c4cdb68577d1f1483",
      x"081ce90cd1d2f1317528c59afbcef8bb157e81b43bbe17d4a4edf71243b269a1",
      x"0e5351ff04dd8a079666c099f4467449d61cea77b65e9c5a850fbc6719ad0c11"
    ),
    (
      x"97d997ff2915ad042c375ce47e074bf666f842c837a7df508d6ef576acf75192",
      x"9312d7988495263244a04315d8bd2b3ec1bb4cbbf30d9345a5bbef488a679839",
      x"9444bc46294ee91ed1140a0f1404a3d7a3a633215ccf0a06f9566429c613744f",
      x"2b54cb4a1fbb0d102ecd6be5e2382e0e1f8e9b277d87b5cbf1a3e5361ca1a952",
      x"41cba8d63149e8d7b3900ab514ebedd53e197d857991cb5d1750b16576400402",
      x"5132fef65a915ce0992e766895ca548843691dce309a4b398e2e689f8dc2f6fa",
      x"82c88cf090590873d41bfc442159fa445e8458fc909192804d397e0937b8bfb2",
      x"141a2d218e283c3cecb12542c8e11f01dedd687419f2a96f8a9cf67943d9c75f",
      x"e2ba80e7d83765c0c27891e5cc76d4966ae44a3f3409e2404f88a1839dd60147",
      x"0289bf85e3a46cc525e36e0923a95074c9e3b1bed6ad335ddcc8d7e7674ee714",
      x"a5711be12982a6ce18014d9bf75b0bc3e87d6aa23c5236af961b616a8b9a4663",
      x"6e11767c4eb5da2ff26935f8e9bbc913692163a3ffdfea7829b975545dc26a07",
      x"212f67c4be2fc59a55fb9c3411ac3e5259d10ac7862653c44cb6f9353e71466f",
      x"17fd0eea0bd8f362309d404ce9f13a80a21842a473b59d5d1eae7f3013bcb695",
      x"da4326721bb310f15ca3e0cde75af6f3c9a02598673cbea9c357bad2175b0169",
      x"ceb7a87c924aa8c9b10798abaec2cb5d490381a35487413f303d4a50a63ace2e",
      x"ba54d1a05c60a36abdcd3419f73aee45910f0565132b8e48edd792f0346dde63",
      x"56bc188644ef80475099d4af83a6b7ed2edb5e7d38e3bc0700dbb13eb46533a8",
      x"2f07106c4bc91324481083e492a8704ed4be1599ca968eab3dc5e87b74ae208e",
      x"cb47ed0db2f61161bb73f9531cf21d33e563a84ed054af93868b23ee89accac9",
      x"c5aaf81e040279cb30495c015d9b65254e187ad02776d9521871de9d25154c3d",
      x"12ecce31d116ea57c52711b369d14d88c721145d609a00f5545f8c858fd8d3fa",
      x"f56220025d38a38ce084a536b386653fd889eec25f9fda7452a6b229733b4641",
      x"b26d4deb7e162602ed1ffe1a417da22a8f17e73d663c08f1bfc82edbd65e4569",
      x"2af95be46e5368f61458074cb854129ea22d839efc5a134691231065978986e3",
      x"0fbe8605a0c5c447930592842532aae79716ee6d2d9dcb4e40acd0e257293a43",
      x"16a1d8d448484965c0ed9d037086488eeb8fcaf50799da6ad3906cd9e0d406db",
      x"9f0b30dd3f0a3f84cb8ce1c887842994c117acbe04c5584b1bc5759583008f31",
      x"1c269ca9c48c2a6720e3400aed686ae800ecbc7e770ce13df498e16895ceb2e2",
      x"dc4017ad4e42d304a965b38f4712778d44fa173a088cded19748ecc35c50e4d8"
    )
  );

  constant C0 : std_logic_vector(N - 1 downto 0) := (
      x"00000000809d4042d802e401d2796754c2f342290e3d7ea97c1b282f0dc8646b"
  );

  constant CONSTANTS : T_RS_MATRIX := (
      "110101001110001101010000111011",
      "100110101110111000000000100011",
      "011010001110110001110010001100",
      "011010100000101110000111110011",
      "100101010011010010101001100001",
      "000011011010011110001010111011",
      "001000000000100001001000001010",
      "100010111010100011111111010101",
      "111011010010000110100001100100",
      "100100011111001000100110111010",
      "011100000110010001000000000001",
      "100011111100010101111000000110",
      "100010101000001011000101001110",
      "100000100010100010000101100011",
      "101101011100111100010101000000",
      "000001000111000111001001101111",
      "011001100001010110011001000100",
      "011101011010010101000101011110",
      "100000000000001110111100100001",
      "111011101010000010000000000101",
      "110000001101001011001101100000",
      "100010000010001111111111111000",
      "010100000000010111100000101000",
      "000101000010100100000111111000",
      "110010101011011000110000001001",
      "011000111011011100111001101101",
      "101111011110100010001011001001",
      "111010011101100001100111010011",
      "011110100010000001111110010010",
      "010011011100010111100001101110",
      "000001110011110110001111010001",
      "100010011001110101001011001110",
      "101000101001101000010110010001",
      "000100101011000000010010101010",
      "011001111000101000101001011010",
      "101001010110101001110101000001",
      "101100100010110100111000011100",
      "101111100110011101010001011001"
  );

  constant LMATRIX : T_LMATRIX := (
    (
      x"3bd7c21f9a733b5860204706180795e2fb9a4262ed33b5149e4086c576778500",
      x"2b1f724b10c1168bf6a08ca9a6226db0229805dd4094b071441ceef4bac34c73",
      x"c2f1810cdc9b2a2b432f44a44439e6f51bb912c0010759a093c504c199ddce5c",
      x"04b85bfda5c0edcb1e479ce570a205686e54c5852ca5ef14a2f95c19caf597b6",
      x"5dc7f9e037f1e56002b2afd28210821c018974358492f3e30526d6b3f1864407",
      x"70ac4778c71be03b7af72af7abb23b574b14a7dfa23bb91e5342b5ba834a3716",
      x"cfcfdb881c9013e6cb0d4db59171b89fad6e6845ce9e5e4b359de8d6328f1f39",
      x"71b9614553889bd792f8d624bbb09ba5ce6be93ec516e53f4245a7fc3783637f",
      x"c40bfe9ca9b8a819bf7fa3f21df366125e15e98991566a12608e61bb46a57d47",
      x"bea8acdde05fad1b1265cc149cc71d81e1bda98850b35c64fe2615ae46fe5589",
      x"6643ff9cd6a035f7e7e2f86af0651d9e95fa3f1b8b24ff6078031de0cc582725",
      x"7059a217f642284c0b7700521063fbc41a6b62c8ad81c9e5f5790a5e734af766",
      x"e629fd005aa8c37c9ff55763289275c58ee2dae904b50468227dbef07b78606d",
      x"7f35531617ed90d9c0e8b3d228a073752e331eec31553d4f3b6cdde2ee7abc9b",
      x"72054be45e615289553919b6e9542ea2c2c93d5ad3f5f6202407c4a8a258f076",
      x"96338709b3a0d325bd25e3afeaaa0cc5afeede0b7e4527066650c392d4a46757",
      x"c3a8ca9ffcd6876760a10c7fd35a6a38eebc11614607dfbef5604cce78046624",
      x"52b903b2fc4b7e08b148a6afb7e651ee267955708693ee225025997aeef73ea2",
      x"abcf564dc7603fe205f16d0e900a9f4d390dbffa7d3031e5510e5636557b97e5",
      x"a4a90e5353ed5792a821bf1301b03c8fba5ae7a2b629d55c97f215ff4f11094f",
      x"2786fc16a86be2ee996d2d8b0b7161959bfa02da911c0d409a946e75fd703cf5",
      x"25a5da8abebde3ba762e76bea633932b507fa230425d9341871f4bcdca06c49f",
      x"e336d4e37457d691faee794aec0a4387372d8f41fd94e8862ce5427722ba4508",
      x"abb9a6a7620957486d742b870d15d611eb723bd0c85e120260a4e927830ac91d",
      x"b8e2af4b00a295f755b700c36fd840aa9a392259585e5c61dc5b7fd4ba189488",
      x"bc6fd5eb2e676b2d3e675d0e0026a4511ac493c1b8bc14b3dbcb254537ea4bd8",
      x"52db02df9543a5363df2b5bada72e7243d4a344be9a53c5c5b354d24800a450d",
      x"2ef4c1be9ff9571d784b5ab1dfe32b134a0aed9b0bb8dd5d521f37ba397a607f",
      x"81cd3e85d3b17dda405bc402ab3c5ea920a160b7656883e402b2d8667bf71fee",
      x"9e33215f545d970d5ec0871027ecd52c718cbc5da20af2e0c0bf11740c7d432f",
      x"583c3fdbdeca95605fd2c21345e1e221b62914f67c45f865cafba4ca5aa62760",
      x"592eca5287e120f13bcaf5676ac7d4a49b4bbf1557d09676a0bba8bd13410b3d",
      x"0db01480949fd450383c9a9988cb69f33d5a16af92192737144eba9af3d3c42e",
      x"2ce7af4c7640c42d8ac3f86e8debd0ace7a1524806d09ed504b75770b02fdcfc",
      x"9db62a5dccd3b6c5c62146ba9dab83d5a415aec40f53b0b0a50f8f6a584a9958",
      x"4601107124a74ac419132ed441de59c9a4a5275e0cde8327322cbc9206395c42",
      x"c70e3d25e88a5dda896e4792e2c6c33aad7468e01e8c5e576a7d8bb9e60755b9",
      x"ae114bac871ace9aef836d843d90b7c024c01f6cce2aec441a72ffe305d8495c",
      x"39570ee0b3780bed8ab5a90a9bbcfd27a52a9640cccc8162382d615c2b0cdc1c",
      x"c75467f40a68070cb413cc74d47635b3e79f42469caf7a36974c945c64f5d57b",
      x"f910da3be720afc49dda5c7ffa4bb29c22e315be834ee4145134fa8da6e6b448",
      x"5fc61a8fc844898ead5e454a9619c34ea040b13c00e5a8e7a116647b87143508",
      x"7755c75eb3f8fd3bc464aabfd869c438870c79710cc535cf0fe80f93b61ee459",
      x"961b311b968c1adca3786795841e73bca15dd8bd08ba2e1e063b47c5b18b7bcb",
      x"3c28104185d43e8746a900cb7b6e61f9dd4027b9fb486f39d4ca2b35ad410aac",
      x"3f859720418bbf0a3061440e44efafd84c6ccbce4d15864e0302465771f89ada",
      x"49c91a1ca58fdde296c11aac4abfd2644fb647611ca7d904319956685f8a7730",
      x"8fe8364800e9efc5d8a7d3ab5cc996af4ad6bd146b43bec3a960b23284f2e0c5",
      x"f2933a4f85601a86e0d14d6b164a2a6a4726dafa7e6b5434a94ef99421a1aa99",
      x"9e42c2568f5791175db2986c960be7563d9757cb9d3d02398f625879bf919b13",
      x"c4e4fcf4391e4ee4e02419f990a3b0877e4c5b40a60c6127ee6ae99eb69b3ae7",
      x"bd58f3ef11c468b6a762ce131560fb7eba93f90f62e3f428fff9fc279d2ba7ce",
      x"712bd13117d36b6a0e77f15efbc3320c3cc9841bd0bd5299b9b6f035035a290f",
      x"e339919edf6b40c177feebe803da1e70f37bc4a1fce1539d18d680fe502b8bec",
      x"3fa740cf6fc9123128992e50b0445a8f032c19186b16c4b84021106ff1c23a64",
      x"20c680d8bac06ed26a1325200f8f29af9c7d4891b36275a86cf021fe1d7fefcd",
      x"b8e8219e870e35fa13d0e95342690b6a489dcb8f7e7221045b80c59e227736d4",
      x"ebbdc5794da5eb5d3b489f24975d544dda178bbdb9684e5ca82f6b4988e14d3b",
      x"99df2e44411ccc1f577d844af3e7f0f05da20f9bf92eb6694a923c2934d13f91",
      x"4127d64130133454f1ca0467764171e5851bc4b62d6640fb145055eeaeecba99",
      x"9b09dd1af9d2bf0c7addac4fe5f8ae550a1380f3e1bda9b387898d2afc7c8cbc",
      x"459fff15be041f3a93cf2aa0d63c45063fd1599af63e5a7bb1eb29928828d49b",
      x"b86bccd46e6749c7c04347e3dcfc05d05c833de847ed181d66e826d47932c4f2",
      x"2f251c9563e584f3b0782cac166c9000f72395b51ec7490308ed7f8f609972f5",
      x"5020fec16839f5e8e2c01b92917025891826cd3d068c419d5069dc36307831a0",
      x"1fc6f9775f13ff0bbdf909fdbb31e424e271d2dd9a73c0e9e2607bbe5c64481c",
      x"cf72d29fa3285e0a964f765dba2280ca2615a30ccb7b0ef25e56e2d561f8e778",
      x"06e615ee7e7dab12ceb0ea948a9a2b4ad4b2e780b88ad36cc80a7a9977fed01b",
      x"92078b88e7f3a730ef487f42737be5d99b794ac2688e70fe88dc2524167d58ce",
      x"63e903b4f284ed9fd7d76a31c4afb43694bbc894835571c73d98bf8dbdbb65aa",
      x"fd57fd3d73ba46f43fd4d34466922a62714e7f2d347d077b2e84241d01de39a5",
      x"f8e7f4918c3f0b49ec881afccb733f14267fa6d6d96932b71979e25aef2b33e7",
      x"c45dfd0c248e2cf0e1d930834fb54f6633299771a17166125879b5fa2c795943",
      x"b713e0866c60fab63a85549abd0ce508a54168a4d3d3fa3cf0381bdb2be15af0",
      x"c2340626d40d5e51b978c16792eb522afda469d5f765986dec2a39c35ea0435a",
      x"4541a58e95829700f309c78b75ac1cda0795fa5b1829745743f1c27fa7236516",
      x"34552e9cfc091f6bec10dc0ed564f5b4a4a66242d463533431b054401264f2bd",
      x"d74a8ef0bd1eae073c011c1d53646d309d9b6a2949329d44a1914d7516ff1cc1",
      x"0e8f8479455eaf8a12ce9e36942f63e2c0824499d2527f25d59f80f2d4c5a143",
      x"46cd26e0d032b016f15ab41f811f0a260e51a71a336076ca4a6e61cfca35fb30",
      x"98c6473ad53306c21e259d695badb8bf3d2ac89f078906a685a7368861fe8806",
      x"41499310ff3c14a117c183e04d4b06a116b01eb5d7123da4cd1947b109518f58",
      x"4f970204b7bb5178f73e5a5765bff9500060c6d1a42e9ecc35d75a3f9bc9d685",
      x"989a6235b7906b289ecadff87d7339dee98f56bac7db9e576fde470ace249ffa",
      x"010314bb4f86474212610d7ee31f557cca883fd984132b756d753df643316237",
      x"92771b84c3b3adbafab84e0ca010f81ddd4fc547b6d5b78ef6f871a57bc3fb9f",
      x"5520614e2ab1c6f943a28dcfa2cac2c33e55ffb2df889b57107efa94a6c229f7",
      x"a969d02f2bea6f9e03fd414bc9519b5df8e048c9da81ed5958b92794956b3832",
      x"fbbd449e4ec2e0f9e8979296f4a508522beacd8f6b49a78cf75b58211b1be791",
      x"157a6271eb27a087b370252300aea24c6df70b3511d3512b9a791affec45c228",
      x"01d0d9b3f74e89a40cff1bde20a6f3e464f0a107c4fa3d0c5db62c347adce273",
      x"c1949aa09e89870b415a8b6489c453176af369e8d0b56df118d4f5378acf634b",
      x"4e2354dd73ea97b7b0f90e9f65e95536fba8bd21f9e64b155015f8707f6f6fcf",
      x"19ec7555ecdbff2ee8ec8c502dfa2798eeef1e7228a05a6c78f4e48837a1b2b5",
      x"cb2acad84d321ba9d5ce98b1de722eec493a63b1a51989ece558e032e4cc18d7",
      x"9b025f80d01584deca2939a6eef24d372da101f3037b839893d1a3b0c34f5575",
      x"c4d16214c336507811bbfdae84771f59b8522738a2633d4ac486bcfb14e272a6",
      x"628a29601d28c33d3196df753b2c449b5b9a793da12e9592ebd9f578d158bc18",
      x"bfdd8411283b9d9f8dc3638c3a432af9a5ab13f175dfbe3b82acad1575bce4b0",
      x"b6bf58f4874ee1cfaff1475c63efd6fc945702f15a69504412c4f7b10d6be4e8",
      x"749a87b9fccf4b80bbeed6ee1c674803c17f392d0f092ebe999556f08973a3b8",
      x"7f6fff9343b55e253bf9cdc232ea0ce4928ef1b827740f37595bce08970ed540",
      x"d02d5c2faa3c00a5f6d8b7d847ddbf00cfcda06655636c515013647372e6a8e8",
      x"65073b6ff7872e0aeb6f4ad7ca5cc5413bbe9cd29ab918a873e754f8483b8136",
      x"eb6d8f2590e6cd739dd51744360d58dd41217e9b2405a6dfd4b1ea8411071ddb",
      x"076e796033d4a4af62248c2aaaa33cc3dbcb8b46c9b4ac78e1d903f3966655e6",
      x"a1bb9fb424246e610e9c3c71146b7399760cb43a734647ee52f540c770715e76",
      x"66db6f214209e55d46e866f5775da4d35d513650408bb729473d23bc1656871b",
      x"591e3772c43e724e42b9d72ba4fa05c77d93c979d3217e868e7dcd096951a37d",
      x"dcf479d2a4f836c819f0759c33e2ed8104a336add1a9b98fdf2d18fbea07bbef",
      x"f3fc99b39c69302c3988c2f964ad929ee98f8f1083b22c677143c66263a47349",
      x"0c455e3ae4449fccaf90e8b5af78524813766a96b01fe9bf8b29248153abd12d",
      x"b5558d6510d8d89a8baac94b612c09190382de6f07bfb00822e0e2a47c6de9d1",
      x"1e8d327a7355547865748e2eeff3c5b04a13d4f530dab89a80ecf3e3d5b76316",
      x"5e837e89d3e0ccd6fe48cbeea813d5ca7120a6f70de299823b02bc73651f8608",
      x"296b69eee876174a3e41431c0e791f30d9265efb410c261c5a36991968659197",
      x"dc2014352c38f6bc96e627615459c030b85ace62d0a86c6b8eb76b935c94311e",
      x"d178cc4cbe960f491ec3792f42ab933959ef42d8f978de24dc3808dacbefc07b",
      x"cc5c2d01a8ca90f699ea0f29566709c69b562d04e72c3fe3238e72c53d581096",
      x"305eb0e7aa61251e63a4a00c93ae9f5d6ae16a7f511c58b6cb4ff8683ae4c574",
      x"34e0c5e076b52f6c265a15de2fa3d621b19ece20497210a666a4c2b6eef7031b",
      x"01512df6ecd5471821a8b38c288941b70f69ae92b89902f0dee22a2dd5ebdee1",
      x"75641a96d0626d8fe30d928c9ac2b00dee2c082dc91eb978165e82737c8e5340",
      x"cd59e76648488d897501d8a281dd55f2659b9055e6fb27bea41a995ba75764c4",
      x"db54c702c469612ce5ed019e780f02f611c5187bb9d2fa9b809e0eb1d90bb027",
      x"0d7319867b25666af41593b6819fb699e3a69a12d3f8616d115166f3a038a097",
      x"e52ccad214623c6e2d682c78f2f1cd40b6fd486ac71a88d1da62b7c9acdeb24d",
      x"8f9a36517219dc9b39452753973f3fc51955b98785254c84355b9ce817c4f093",
      x"0034f50ef87832f25cc6fcf1dff0aea0cfafb26ba789d1e082361cbd4d0852da",
      x"bd9ab431280a02c4ebea15abf335d8018d25f2a98085f192a410099e6f1246f8",
      x"e1ef0959fe4fa117e5f770738d560b01929928c8bf5dd16662d90e0ec9b22866",
      x"4be46231a80e5df942cdfe1bc33a94883cf80f5bdde869db681f9510318fe8ac",
      x"c446c223751b971804977866ccfdb2d59aef91e9d0bc3618a2602e6d14dd8723",
      x"80346ccd9ce8f54465a928ccc800febaf5c5a08e7190e3cc3c42f8f0839af37e",
      x"4625721633cde2419ff34f4545b8a3ff8779071435cc472c66537505256bbf92",
      x"837a1a16b16db58b418513567e56f92b68e8aae4e0d1ab88e4256b5ca019017e",
      x"22b5e2772ac112273de1fd80b30952844cd5b2b905c053a4b2ad4d4f945c9112",
      x"2696de97d9a609231fe6a827272fc4694a784a1d400ba30c3adf83a1bda9bd78",
      x"c9ee882b04bf09cce039e1d97decf2f05c7379244426f1dd6e7c59adc5f74696",
      x"11f7cf0085e0e616d50b1d8d70a1139af6fc9188f0898857564fdb03d3e6d539",
      x"150e0ddfeca74b5f979d307c563521e7af42d4bc717153576994b452f3eb613a",
      x"43cdcb00e0b91e936110212eeeafe4b7239caba64c029353596c7123130f1ae5",
      x"8cca09177c924bd1006b4b7142e4c06118ada80829b50e92bac3f29fbf8fe3b4",
      x"de21c9ae669c7b7167c8a2452b9d960c5e0c27ad1bc86478661853b763fa3769",
      x"362c940937c94e8a159d09c18dd0822c7a8b76fd4dc450de54b298314d329926",
      x"b27a7e18b8e60add0cef3a2a289997a00fb01411a316e3cf0692cfade6e419f1",
      x"e3d5f465ce229791106f1d2d45db06ea33237793e38ca07d86744e1678e6f91e",
      x"d83df49d065337fc144ffd2a91a9c1570413807a2e9865621c3260cf531c203d",
      x"d4b6735668e268aaa131deee5758b434152c372728d788b4400d6d0fc1b8ab0f",
      x"52e313c5240d33a95a9825505f67d7acd4bcdb2dd9e9e7ee089885d2515104e0",
      x"eee382f9bd248d7baddc8b0a35d38e3b58a16eea0eab9375c1dab5eb826dc6ec",
      x"c8aae666c932f8f12e31d0c4b088e87d693ede1c107756b5fec0202f3a25c052",
      x"33764f63e7fc07c87b1bb68e1f21b63fbe4455567816da21b8739c1d1c2ff033",
      x"46f28d802b28fbde6c9cb972e5b2353ae8c65396738ed60eca2bc8fed8e879cc",
      x"252e863ecdf3195d15436d4afd578353b7bbb47a8d03f66d8942f859554c96ab",
      x"8a6161b75c6c32c1178907333c4097f113f9049d21a5ee753acf31ff1db86288",
      x"6eb54cd0fe8b2e9cee9bbd21bf49cce2e4e1633908747464b8a6120f08793a0d",
      x"df2e59af2ca9b1dab80175163c0a5e06887366b9abe16f9128bc0a77774140e8",
      x"5b38a874a90d50e2dc06860a98830f6b05cf68c6d6d251462ae5d0ea88585e4e",
      x"636ff7f1dd4bc9c2620c5e840a57109093464e601f0a2c6c3d7d246623649866",
      x"d6ef40e755f91ef207c356107b1bc0cd40f7069983a6453f620e5e17216a2ea3",
      x"9af89ae1ad95af450acb8284953de5b6aaf59efd51bafd29e004fd559029d003",
      x"c7d643db04ddf1b32d618bf0ab6c2169d6850b979b0ed4923735678921ed1c00",
      x"3b99a10bd8c53ac4d237f32cfb2f784ce2d7a48c5b67746115911009aff706cb",
      x"1a8da57f27a7f5ca823394a85a3bf1905869f4a847a9df808283e73d3af0c6b5",
      x"b5863b15acf8f9856726c4c3153ffb9568879c36db796b85e159d8d420762b29",
      x"9f86c9094f0ff35a60f16ddb4d9414693514c11bc6bcc9e6134cdd801bbd841f",
      x"4c310ffde836e805b092b937296fab0087eae5a3ba1d49326c2f6477794ee529",
      x"3b6af05ce1673ca0f6ca14e3c41a7c0bb500faee7829fba147ac80d580597c93",
      x"4460f59f7cc0cb7e6453c4c2d200d0cba552d056368a1919927f196c3e322bce",
      x"1a3b5c943a2bd6595b10b52a24ba1c25031ad3ee19d4fa107b52ef9a21f6b1ac",
      x"b24aa365c6c0eeb067dfa6c42ded065ed68714b0b47a586361d7da0d12a2ca8a",
      x"7a63b3a21d27a0300a53a5bd7c52c94fe1dcf43d303e20e9734136aaa5957837",
      x"3caff05d8e9e999b5e06c47f2d1dbd33ae354fb21f0efb4ed6a36374c2c836e4",
      x"761b3988f70aad175d9345f4c6e3ac9f19d2e8c3a2d76d01614e72f4ba4fc97b",
      x"47f63c2ca12cfbaac9ffbf0a5e26f552136e58a74ab6dbab45c0ded253a1b9fc",
      x"1b90a07d68ad18354d2ae538996f91be23df74260714764ac28b7cbbaa0e8713",
      x"a63d99dedaa540aabc4c2b8743dffeb1f161866dc55223431fd1dea6f8d6db24",
      x"84500195f5b7218f4d3a677a3bae2ef1c9260cc848196473797f6d06284c2e4b",
      x"c89dbe75c698d2b3e8aa73e3830b326484dcb0cf982b9148812d73ff43377115",
      x"a21dad88aed51b44a2247fd64ed60107a24cad5852e5fb37ae5ad66f90018f8a",
      x"e2f874fc0b6291436e352006c33e9f0e9312dd81cb64c850aafa43de69a1ec5d",
      x"197cb4e9e6fa2d2f47ef101d8a087d6a388d9e9a66731e24ceafb2ea6d38d9d3",
      x"f4035d0f8f65be5ba7420c7a07efd9c67527ff9e15ba40d1bbdd98c88fb13502",
      x"12f9b307217b42f3cbe2220fd2d3229dace224dafe58cdb4fa15cf248df7bf6f",
      x"4a09fe4afcb4a2266c0aad2acfdf2c5e3b54a1fe2a0e0e691f511b7acae3a0ec",
      x"2132f5025fb0c17e5ffdf6b618b5c40a53c29f96981dd113b1fc99cbc779e398",
      x"90b348cdd194ee1308a68813af58ead387961a1c50001fc50719ae2e61191b4d",
      x"35a2996693bf5df6bbd00d789bdc56eeccc840fdd007d771b61ec733930c817d",
      x"0aa108b9e981eaa3c2178841b65ffc7646c5381f445b89673cc1abaa4df78498",
      x"2d621965cdb2fb550417e6875da60ce8ea5f83fc2eb7d2969cccc2d200a0ff4a",
      x"52d47a6adbcd915cb18cef09cdfab372387aaf09d63ffb8b8027f19e5f15a3cc",
      x"9dc443055c2a20f9a1a78db042208c777edff40e771a1c0fefbcf9fab943215c",
      x"4bd76b0374597bb282f4effd4fcf3263475953a24881628d4f7a20aecd24c35b",
      x"5b0b6703b07d41089a0a78d73ef85a7f68540c16b1eb3dba922460d5365c786f",
      x"c3cffe93d065cdba36b9b72f2910a8fd80d5b9d1244a86d5a760c05a2f27669d",
      x"0dc852abc16f0e0670b5eba5bc6e7e0e7a9dd09f7fe9afb3b5807ea33a9d29d6",
      x"1fb4765e70428733753f85dd82d09070c8029f4b18a6135fd5f6d6754707b533",
      x"34d275ad8177f2631a2d05f84125593d45f3e7b78077436ce84f047bb2053357",
      x"6345563101ced7b113cf2abed5cdf13e794aadf410c8b6743125886b0a6cc78b",
      x"b8f84daae24fb3ee2d6ce870c9cd91af2fce168bc4d7059fb48956186be8a39d",
      x"bbae7cd662d0f799958afbd0db5aa17766ae2fbd975fa0a84daa250582bd760e",
      x"e3f2076c0c7f9ddbe98067617b80cca0d9545b7563ed08a45bd7b2ca7aa8c3df",
      x"aeb47014d61f67b1937324d3adf679901aaceb2a4bb739f029617a8d5a2d494d",
      x"e11f07294606b4a26a36cf5162fe45a466f10f16f1cdb19ee243ff78a1c3c6fe",
      x"411a3a4e4b9fecfec194b4ed6df9ad639afeb0f3ddb27e213941bfc5c06a6ffc",
      x"8af41ad088c76a67b141fd7b4306a71618140a8ed1f1ff10c8a27a374681b26a",
      x"72077144c22f4df448c7ae19b9452ece7e18a0e7760f1dbb413e7d50f4031e49",
      x"ad4083e4df4e67a7aaaaf1814b02d1565fe282e7bcb869e556d2c6bdf41843d5",
      x"e2f8f46eee43c9c88bcd2e201e6d1f053023f3fad23b11f80308dd205a39f1e4",
      x"8d2c24168b199237d268166581d03c8b045e5d47688a8436c01b81f94cfdef12",
      x"50ee61f98b763c5badb1377c0aa969c7e4a6c1722ffc7f9eda142978252d70f3",
      x"63b44654cbbf2b877a9df7ea5c29712be76d037a39d95efd09e26bffa82334ca",
      x"ee22a027ce2c49f61589e6feb1dc56912c860cdb51b78bc6f52061ca0e40563d",
      x"8e4bd10ef4a5ed511a76d4006aa70655debc38d685c83641ccb476c016f7b860",
      x"3a68081d1f75a1bc2587dfe61d9aaa14729531e8dc2b03b69136c82be7c2d2b7",
      x"7a56d539330c85abf3cd47ba35f1f1045913b879e3fceec1223e126504aa847c",
      x"ef8d4bfa1f9cb43ffa1729cc326911bc4778cbdec320bab4782859c09aa5abf6",
      x"2aa92c26cf58bf25d7a83458f14168ca4f2cd5189481b54f0f4495836da64b4f",
      x"1d3dbdce7d5cf65c21adaeeed527618402835e8671c280593d1781e29187344f",
      x"e3ab4ef238d8bdf2eac498a200534a0ff891542f509e8fc2dca45be858984966",
      x"283d4dbe48ccafa16d7ce4d163e5221e4ef6e660bb7a6ddcb9c74f789038fb0d",
      x"00dd35546d5204d1443d3e787cb574b9737c550f0f6f16370f3f5350a06cea90",
      x"a921a507b9f8e0f47cbb30641bdb9d88bea22474b2388c2826ee8a381cf18ad5",
      x"9f24490a292b40410820341eab4c2ebb469c2f967e237ea4d8a9371cbae7129a",
      x"39e0758660efa7e3577e40f645138326911ce45b6806c6994d96a716e6d18b2f",
      x"8fcbf4e74311f40584e7352efb1803248c1959ca9247a9d07bf21d841e2cd20c",
      x"8a62542f624ea545ed178a5f19af246293f837828edd15621684036753a614de",
      x"1499c8a9bd7e8867545e3183072c06086dc5a32e1f793a4b8deef43b9189e3a4",
      x"aa8992983f7428e59cbd310a0e74d7a1575d31e568831b7dd245071e46124962",
      x"24d90d3935635cf5881c85e08a6cf0cbf3c09b4138874c754803b9b7ec877482",
      x"28d1753fb75ea8ce976ea4f3ab65b3fa274e79d08ca4e1f7c205ce02819684a0",
      x"78f6a113f21142b1d43d2351667fd79e5fa8428dff32b0f87f5011d5a7269cac",
      x"6e581f8e8eda4823db3769d57f50d2e2ccb8d00d36000c3d1abad444c3389874",
      x"f10a0519de2bb2d4ea1f711691c6e3df856f0238439084fa0000bb8193ab5be5",
      x"6c873e4ddbf416e41583987dc6fedf2802ee3b782071aa102025c4671ed40298",
      x"e57f12b6845345c3632713d0e2f09dee959e199641658a2ad94375610aa29b74",
      x"abbf0e5b49f2d4be436a101d748433ce5c5fdf8ebc7c327575d901dac50d4f53",
      x"16a7a5a8d3fc75b7d72932cf10dd6a63581ee6827979cc62620f5637714c2c6c",
      x"1522ff0b7320fda9b7c12e5103673a6cd378edd27cb69131ae157ee4826d8848",
      x"b6c714e154b4378237fb03e572dbe0b380c2cf36dea3ac37e3f62464a39c6028",
      x"3ab029c2158e156f7f63b0ed493352a3df6c35705ab4f3dd8c42d5b880a48ecb",
      x"7114b151813490b006de8c7b3f34dc7626bba7771c407a695db27bceb1bb11c3",
      x"2f0f2d86ef8b443855d630fab75ee77b7e10d1aa87d12e04313ba37e29c6190f",
      x"a8ce387c51a91bb2c4a0330607ba0e30d30486f502d5f8c52006b4f3084f57de",
      x"1f61e762f1896771926ce0dc0118c97fcd976d276642f7e8a7f3a83b15968e03",
      x"01c3929d693145db2da6a9bc6457a49af4113301084c595b1cd92d1d62195845",
      x"6e34dd4cd1a970db5c4950a3797702e220f65ec2b3e91429f6f78a263a89edd7",
      x"01618ce073aca3dd3c256801c67022f61b26e33405dff60b52b559f1b9857d9f",
      x"e1c69ec27020a9ccbc6bb736aa73de89b9ff59ae92809ac82781b68b070a6c19",
      x"f4b73573261a4ea79b66e85352966bb817fe252fecf594aa952b38b36dc454b4",
      x"c10ce703eac3720a23df1129b8e84383d2c79c3e69da0ae4888b78b655197710",
      x"910d34a9a1511f64ff53657787038481f79dfbe62f5929a5ad79d858b022ede4",
      x"69e052323f4380e3e92a65d0359d95df73c8bbaee4a74d8bc41523bf353ea55d",
      x"ed444206d485ff14508c8c8f1eed4f2671667e2b6c44541b38c415ba69605686",
      x"4b056980cd707ace501276029d7320d0ae452083a456d93dfd3d5044dec394a3"
    ),
    (
      x"b5701ce140e831e5750344991c260addcd0fece2dcbb0db48371438ba5455a33",
      x"7c170620c84ad1eafa168c0298de652bde3d338e0d324847e4f5b0b980ed677a",
      x"a4242445accd55d9750b9cc13cdd9cc0827a528af7780c919e99bd3f60ff7399",
      x"ccfd99d8d14a296040736b439bb7233cac27d5c7471b194feec5824f08cd8f03",
      x"7beb453b9b8c6ed91ac8a4f3d58fddcb762b426a2de91791eb6b99f5f9babc2a",
      x"51941403e50e169abd742347bc7f3ee6fb974d9bd7030471582f8266f7fcf129",
      x"7b23923e49f6cbb4de311e67f2cd748bd45339a6a0df6e4f62f80acd6fefc48e",
      x"565ea209b1dee40d19c2ab390730d5fb4a8bc5cc75a0ba44985b505ed03eee96",
      x"3e010b0d7c990a7f7a2daf512dda264edef15401af23ea824f1c7c063ee611a9",
      x"13854fb5df43d1584350244c60ed5f32255249fe762424a10634c7be814c626c",
      x"1363640bff1ad83bc3baee7952686b4af79f44a5d361e76656a9f813a93d74bd",
      x"d8f804fa48c706324387adba4aa3dbcc16b5b9a6c766011b3068ceac2a19436c",
      x"2db423e106be571bc42ca02f6e0c565b4e04b0b6da8a3b972d340fe4b68032a9",
      x"0c0f1476709d4f779a14110bca4212dc92996a0b9b77e7f64152d44f4aa7b8c4",
      x"eadf1d5a43bd97c62628760a58196c6f30c85308af2e3f8f7086df42551c1a3e",
      x"22d9adbd53b569d852bee05e838d23c2bd15606305c3cb922273efde6a856baa",
      x"1a4c8f7f657819c5a595a7ddb19c8b5491426cceef1cebf0512205765b8ed258",
      x"8a0af93aa14cbd8da3822feb7deebcc28cc55a8e0413389725cb80668cde7a6f",
      x"c563d6011335356ea15a800e355bb6e6186ee5957a9db6d5917e545c354c8d76",
      x"921ba707f3eca8769ea3a922a5a83409f50feac2249f7ab8f3ae8912267d0906",
      x"c13f900546c428841f6de8dab290805cd5d4aee7489a5c37c9e846fdaf22f1a0",
      x"8cd4867da01608178304b451af76ce8e53121d002c9d53055996a020c9124255",
      x"0fc3d215b2b8bc5b8371391d1110cf7f9bea0fb077862f4c99ff86db74ee5a37",
      x"3ae84a5b0f5cabd6e6ecb6559318448bc54dba559d51d78b2208fcf85609718c",
      x"bc5f1b35155ab1b58cdfcf5398c4542044e2f865a26aacffc3675dcbf4f6c31d",
      x"ece008def686da5c29c172bcdca6979f2db584487bf81ac996e67f2254fe60fe",
      x"9af1da6d844f61239b18fa3b3a7898bc803bb879441ea6b96fb99d706d305ed5",
      x"daccd2ece7e5a95cf57b791ff465355d549969883a2aa58c3f94fd377e82354f",
      x"c3326d8ad434d3f75adc8f3c90c571b823f0c632e7f476868806bcd0f5c5eb8f",
      x"1a378908a3569924bbb59af5be4a07a5ede6d2d6470caf654c6ca69e416ef6b6",
      x"2191de7cf3544fdf89e20d21f32da5f4c155f8fd2379806a4208032dd1487a71",
      x"b6f0212b5b7b5728029a87f7e5eb16dab31c222bd24af63417f0db88e57c3739",
      x"49578831362e4c708ea1320e59b8dae258a3aa7fbe84ee8f91005a03d706c3fd",
      x"7f3667da5ba4edfa9d7b66b1d79583db220a11c17c206f6107c71e2010a0c9ed",
      x"0b367822a5db36da95a2df50128371050d931a5de3faab55999a89d92652fb84",
      x"233e721fe44c5f3b0326cf9fbd57ed2a035697721b7fd06cc299b8736ed8824c",
      x"0c278a9e2247f11ed532be2fee7103bbc56904f5ab03d39cb7108af0c0557236",
      x"f6e8dde66ce0d77b0a939f18a0c94f84c949d15e9edcc85bd5b00af30b5534c6",
      x"7444a7659410c502f318d3cc21dccef0b0c49646eed5ce5e62e0085a5d21090a",
      x"8e5f04109a7229f9b27cf390130db04abd2d17c7c13a167fb2aaf5c02ff391f0",
      x"c3b06068b8268e48cfe3f0f3927204f88cc454e747692a882811fbef205ff368",
      x"741043bf2ddc1a8f1ec79cd80b11f9fab167dd181324d0c7a6bd19349f102c09",
      x"f0de9d1c202fb405414350e7528c7cfb03b5cfad89a2c10b8837219531d06da4",
      x"ae0181a333a60bacbf4ab6e07e010dceeb03ff2198df4313ac594e7c58b7762b",
      x"fa7d17033fe8f95f12d2d24e120498d15ca002aed498949716d7a1f31a0bd78e",
      x"3b5941b6a9f2b1c546e23f461a4eb2c4430274834e6f1b5c85a4d862fb88ab86",
      x"ccb960448b0dfd9d89a620e75f776610ce8cbd1cdca081622db97f30dcfcd96a",
      x"96b10fcae248283c3532c5d78fcea8cc9ef6d2512cf606ece8e6268c2700e56b",
      x"c92af82253cc35114b6de1fb6bf015a7a19a9f2a5917a8c509ec4b2abdc6f59d",
      x"77af852db0452149d47977316dc704e32a0a1df1fd7aa8352e44d27e2e8921f6",
      x"e0bff048b3fe332b831603b3d3d851e0a0dc744f394968dda5a06f1f9339de9a",
      x"f59ca36af60aacacf9b34401ea1cb397e54b8fb337590c4153c8fa48ee075d53",
      x"31c5f4c1b0ec7e959f9ca703cd5e95503e5993be6bbd4b156d22fb4fb345bb06",
      x"4d7223eced6786fa1895900abd7045b0a5d929e2987d732e5e25dedde3d9e808",
      x"01c7bf730cd3587c3005964a6b419aa6dca0707cc44373b98d1f18317cb99675",
      x"8b467dce3c5464e0dffd44f9f2f04415f084fd6c46b660bbd00ec7a4d9750ba3",
      x"650fe3e93acd9ba5774a44b9b7d6d0d6bbaaf27e3f308a8cd9d0c671258b2718",
      x"ec8aee86243213d0db6674b78efa425aad8f76297d15904d21e202443a0c51bd",
      x"5fbfd2326e3b4110aa438557b66d3c06c384b74f5fb8138c1f4a9ad52de4cc13",
      x"51a3e847c8770833eaad9355d0d000191aaad7ada32bfec39e0a45ec3d8896aa",
      x"3efa51f11f7cc40879fa1116d30bb844b8b864ea954ebe5dc9b9b87b676c3529",
      x"68338ce22092561d8cbf0654cefa18a02f3fbf07abde643b3f3b05aa3c9ab091",
      x"687540eb7c13d4d4c2ef9f74322c0d90b82a2fce003dc09cf8ad70e48d422deb",
      x"f58de7d3f1c06ea7832e3fb77cbd6f36cb985c247676c6570ff422d577572688",
      x"91016bb2def0d034c9623426b72850e7be657953ee143ead6903de56736dc758",
      x"7b8d61f591e9ab5d93c4ad5788b85629748c3b1a18bb81d5b46e41c7d4d8c64b",
      x"472af5605bb63f5c916272b06493404844b6e2b29ce8da425fdf8f126e8befec",
      x"d8bb193ca25fa6bf4f5086af31e7d7e2396b2dc95f4ab2c5a4a0e25af571fa7b",
      x"73a689dce6ce5e7a07302f75ca6395cc53d378eccc337e355f04dda9ef8723ae",
      x"84300697e6012734db082dee54cd7f51271a7e5f9290b4b20b9c2f424e0eeab0",
      x"79e61940d7cea38076cd81268cda370f2adff4556deaf4b30f6c24f3e27e83c7",
      x"690caec67085d25b89e56344586ea59e60f31197f38d12eeacbbca2d037123db",
      x"af199726691a8989279a5e724e5cd543c73efbb7df36b7e3282ef564977c2d54",
      x"56ffa7e7ebabf5654011aa991ea47f7500c69c423253a7d01863897f2f12e1a0",
      x"f8b1d8ee7c0fb7e675fbc718402c09e16cf8e0832226368fc414c70c4e3dceac",
      x"0adebc064339256a19604b4f42c6dd2c8adf8eae686e026a5b48c9a642af4e15",
      x"e8167b788bd7ec58df47d4eb3dd418ddedbff874c6d94a3ee74b64f84164aac8",
      x"acaf3473c4ed249c8891357cb63bc54cfaea68cc3486ab45a8ff341d64bb451b",
      x"c4c880de81cd78dea85053b2429d20758c8fafeeaf146e9a6ccfbe780c70f215",
      x"f8ecebbed5fba6bdf8476eb711360e2bdd332e47fc51c92b27adb54c0a36d524",
      x"be194b59b0b5ccd167533a2a0bde7ada8aa7771dfdfdba691b2a1ee6d103f5e2",
      x"70605d2e66408896da6b8dc597b3443cce723bc25625718e86fc458b6565018b",
      x"8ad799b40f446d3f9b67d8b8f17275b6233d2295a9d52627c55790ab1289b562",
      x"3fe90c9aaac838c477e95ca45be3c453b909b58830c00242b58e338eb5233af1",
      x"fd28ec8c7e6d5c17c0d35ff7f2bd8d52471dee36e812a8f5f5a26821a68eac16",
      x"c26f9b87ae0e1cdf67534955e8a81b0408bfb05c6603b6aba3b1ae391aa76867",
      x"6371c7f12f73cb42fcdc106bba71d8e2962998098caf0b2e874028a77e50c2e5",
      x"c58d79d58ac11749474ab73b37b9c4eaa3e243e266d1e4a2aad4c4e192c1d908",
      x"d5111ff10846ca94f7553e4d260335dcf49c4f15ecaad7e0f81510a0e3aff494",
      x"8c8b4700af59cadaeb0d2e1815691df362c88b8c12962389ac2d2aef62f5a379",
      x"16f41a2aa06cdaf5551df3e6d7b79529806dcee0b96d29a7e81c5a7fd49df475",
      x"b67764c33829ebd727bdec370d710309587254fcff6bd5c50fb21c8b90c1a626",
      x"96fe74077fbdc11655b2ccd4090617163d0fc7cb70ef9b33e756d982f2e4dc06",
      x"04725bfd2bd900300cc3bfd29aff0dff159f5059d510d567f9cd7acab8cad582",
      x"0b0c4c1fba06d4277ce21b236d07811bd40cf6ba850da9f17115fc62db1352fd",
      x"7426d809fa170c3e4a8c469285cab740920b18032a5f212bc28ea52f1b5482b6",
      x"bdb69958b7232916ebd0082c6608991df38674c7e71d48f8541e8394ba156aa1",
      x"618f7ebba8e673717d9c8cd7f947e1db7dd22b0ab724328fab33e38c3e7da5ff",
      x"4d486ba9eab845f712b7334ec66bcbeafefc22707647c43dbf9b942d8d64d590",
      x"61bc98bfb9aa1d0dd38f2753274ae658a350d0dea4c74cba74ad28ad7799a220",
      x"85de765d72fed374ff29f836081aecb4a5e74d43542a74a9c17cebe1da9a85d7",
      x"447323f91720b7c1e2d67d642a1f683c6fd881d4afd761d14c5760fc0ad0a1a1",
      x"b22ff75918bf0e9846e1939b216b03a3ba36c6b780c38a87fab608238dbc52ce",
      x"ae9a03310fc003cbb3dac53e9e42f479b7559229df430f8c8304a78d7d03f887",
      x"35a06fad973a6fc96fa725f9a574f23786bba07420252cf3c5e790def4dc17ea",
      x"e8470e66e81c0e85bc26114e26bec0c28f2391697693c9c4a4c7a7be12560de5",
      x"fae7a428ef6a92c5b641ecf01bf44f5b036fee51aa92a9bd2fce010fde72524d",
      x"108890b579675ede22cb796d7eca49ccc31200df3ea8f3fe7f787470c2dff737",
      x"2bc62d189b5c561c7d72584a2aec2cf661c32c7b5b615f7eb24c3b1efa491942",
      x"e9bd1ca64c9630dfd4eec835fc0d76180e8ed0ead8030f74c7ac8d485e9f40f5",
      x"61ddb0e6209d332f0562c53f724c3ea6a5c6809f5401193d261775cc764ab767",
      x"a6f5a8c8d41e25147005f60c8f03a918a0006c1129d7747189277a1cf40fea63",
      x"bb83a8da0378bb67dab32d10f58ffd21f123707495667b4c0663b1488e6fd7e1",
      x"a266ce104c5e0c84e2ac2d23df56ee8685449504821e981010e2301ce4bb3d4b",
      x"23a8299de0a92045185d93aca463cca03f65ec6fb01ee73f8e23c0e7c0e7ae0a",
      x"5bd0aff3f8c9ef913dd2580b6e85a5c316afcd0a6e312e9bd32e0d5be2f413b2",
      x"1fa890565326b3a7432aa270a6a1a04222f66cebd91000962c90dd083cb5df9a",
      x"1593330cf769f330cc136b5147a069daa6f0274abd091fab1e9277677906c0e8",
      x"74b4d9448d02922ff8dba2a0992606bf3169a6df667d8a85318b75bc27f3dc9e",
      x"9b903d265d33342add117a17566e91a3885e77446e0cf7a191fa49f04c51feae",
      x"727ae424e299deeee23cea69eb5b6b6d0b79101c796afc7dd97f2a1ca54d6e0f",
      x"766742a67443187efb2e1b946d470ccf57d61b3e1fe00f86f710477d4634b138",
      x"45be4a74997cff262c93bed8ba68c79ff8c56c082dcf44ff3ace5bd9adeb0f46",
      x"fef77441014eb5e801885ec0a8c8848a73b35b91301354edb402df8d23a425f4",
      x"b1e799c4778d57bf2cae80639e11c1381a04c0fc24b59abe13623486e5c53d9b",
      x"a2e6723b0e9676625b148fa481e59f568593d0ace5fcd8fcfc1884afcd08323f",
      x"74f3cad84f62689f2bdfe9163672f0d86cb989fea2d944a7260547554e601f19",
      x"2d952054545c60e95fa90226cfaf02706c5bdc3c795bfbb85ca2b9e8d3e342e0",
      x"57631aa829a4e9a6f1f161d723d551e9eb7ee6682fa55f04e05e07a84a4964e7",
      x"8ed8731527d930c4e0e892fc10010a2b16e91623f5e0a9fa3749cdaf59841aec",
      x"514eb7b3a2997dc466917f70dcdad3ed7da1cc13d47d124c5372381513646210",
      x"48f3dff977b43ccb9f2fa34ef692acd7d82717aa90cddf71f3809f517174ee01",
      x"3dd6e6eb817e83c041da5cafd3cc0fe786d5ff9d68df706babeed5d6b19c1135",
      x"b3bd0fb0d4b3126c9c3b450c085cfa30a4bafc3853cdc1562f843ceb0e59dcb7",
      x"f5955731252e7366eb23820f1c52cd617cecddf0919a0e35cdb22f24e78cc09e",
      x"4f63524833575288ac3f7547f3a86e489360c790415177afc516a960898a527c",
      x"c6c0bb513975d086b9fc0d8a8617f5e9e071617a765ced861894cd488e1a9177",
      x"cfbfa773a53a4b8a025de91d10b485b441e68a8b314c69ae447960aa74b15c50",
      x"a857367d2429715f4b74fb4661e7e0209f9d49172e888b861e6345716d48cb3b",
      x"f35799642ac0e73e30f65319af86863e627da44fd1dea0146fb57a348c95157c",
      x"6840ef5f6c2a8bf6b13dfacc5e02912ef35e22295a37d1536995e6812f0695fe",
      x"6741aa916f13c3c574b8e3628545c0dd7df0ebeb8b497a3b5cd18974db2554ed",
      x"7a89f7c80c5a3f39cad418e28261ebb306ad776af92b0b802ebc44cf2c4e184c",
      x"c7cb5e43e85e097a32ab6d0e0c27309c8f2e8012d25f83c15b453888d11edf9a",
      x"4f31191f014e4845030fd94db7235b970a24aa578a3d7df21a0abf17ef0b8a75",
      x"0b2ea2eac2ae9b76346d31e176f76d7d4643b8088098ebf9978234463d85aad3",
      x"e715ffeebfdb257fda951eb2f45021589f8648bc1ea8222b39f1640d1c78180a",
      x"0ae04e644781a6b2180da8ac226e0829c5f42fbf967cda576b8afaec14a88ea5",
      x"0c9eabe9ea6f12000d20e1c1d183470d18cde22a8be8998ea2edc21e49042a5a",
      x"26c69b79b864964a9f0380788ead3d237016b6df158a74e6d2b1987aeadced94",
      x"16be82ae330946ec4b33ea1732fcf656793bfacf1180b371c5a1726827056736",
      x"ccff7d3c8b3b501897f5072788760fb7640d3bc3ae5ebf30e7e140e1d59c5a66",
      x"29d01c29fcfc7493b64c4bb57256fc5dbe81e4b26aeb1d5400e8294654b015e4",
      x"fbb5e6073b34bc84ebe1df4c27402d7302f958c6d865181f4b580a62dd8fe7a8",
      x"c88f77c0e9ecd8b1a7fe3a5054e3ef01a7fd4e5c5b04a9a9568340334ddabf69",
      x"0f433d642a8d9abb6d7cb48c8b452b953fb40f2b4c7c5d2c6166f39d46f39cba",
      x"1704a4bab1eed061d6f3da9c82a6a435851044b41b438b743e6c4ed841a0c55a",
      x"6c4718069a666e5e458eed78c4f303586bc1f5071e8ef6e9b17e54152c11f957",
      x"c1e025c90a1adbb33ac17dcd7974f0994277c70d6e2385f81524878cfecba6ae",
      x"d3e8dab28c482d54677e974dfdbd67b7be41f57d651330d487ccb9fb17b4d1bf",
      x"4ecbfe54690e166b6c2cca89efeb0828853a36814819863af52de0386a208152",
      x"8d73d8b69674e9ece90b79c915f36eb854acb6e1ae21e37c3e463774c9a7c117",
      x"56be0efda165f89b9a652e15e46033a19311f6fd55f6f16fe180be625c5b6c26",
      x"18f8fc9384fafa6c08f4f3d3f2b3b421092fad38a4d0e0851185d7db0066e61a",
      x"d3b31980e6b6d24dc7ad3dca20484a77516d2313a39bec64f7b2c73bb6ed2c56",
      x"dd626b7099286a3d64ffc1b1f1ede5c9d0644f4ca01c908b78e63f7317103e97",
      x"08b1ff509fe587a64fa6417d2c0fb31cd5273725383156f844c5ce7fcd70bc8b",
      x"f1e47f22997a55f614ee568c0d17ec35a90f9a8383e2fee10e527c9593238064",
      x"0f06dcf62173204577290632250a7cea5011a966ef94afd362146b146f5ab50f",
      x"84cd3731a6ce3ae587acdbdccbbf2d89949fac57ca044ba2beadf4fb09aad582",
      x"20192d5e43bbebeb1908f56db2141a16419e5e192299a71426d769f3fac08f93",
      x"9ca6a80e26040fa3061e41dacf047bb053a1ecbf30e8a7ac29f4c3a8a0c05879",
      x"0a17428002ab80f75b9ddc86a0f1bf386cbf94701abd1256523eb6cbf607a23c",
      x"fe2ec261ae1202d581ec3c3279c90c967defcde9e6b36763aab88da9abc992e3",
      x"653eae9fd56a1728461e87766ffa7efa8a07a23c42eee48deeddf78bedd6d08e",
      x"daaeccd7e5482d21c21f0e239911067b008c0e7b35684fc7ab0712191482a3fd",
      x"e5e9607b08f2fb687354d0191df1ee54e7742536e070dff2ece82b25b7d6264a",
      x"09d8b4ae439c2f51b8c39ec1d36faf63166e12068e973ae7400a0c5d24d680df",
      x"e33d13a8cbb34b637d3eacb5be9f9f8b64e1d5bf15591e86fb65c877e5d3ea01",
      x"65949e4135db4834095c42632ce64d43bc032d3e608f269d98709aedbf54b6c8",
      x"90fd4da47ca0ad06beb438b71fe743d3fa2e23146213593933105c283825a8d8",
      x"d045aca7cc76baff472795088ed186bd1a89b781c60624f6422dba7083ceb91c",
      x"5075302c870c3e46f5fafc25ad00fcc25f33d4c9eeaef5ad4e813b6e3c30f2fb",
      x"008cb931af1e9b5fa547c76797629ef81764a044c1472874a499160c1e74111d",
      x"d74894b16a582e6934d3b8b4c77cd46fb3e534c78fb272e0dbfc713c70ea2435",
      x"8f7ad827227d618735d119d82125dced576108653d649ceef5a12bc3cd0b18ad",
      x"ceb91356c7fb621dd219f89ada27b96263a67f61c37fe24c36c3274d2aff6386",
      x"d4f39095d9b356484cd22cce0120afd6c9381927013bd945187c0364c0bb0613",
      x"a2c65d1ff458f085be4dc58439588d159ac6790b08467973d9590c9c8ab07612",
      x"37124f650eb9bae07e8e68d588a1d0e2c6dfe301b49c686b57629e18a2c95897",
      x"d1d734b38fc2817151efafa8da69b3a385ef764c20750aaec1c7c39023867b4a",
      x"428bac7609c4e652f0c0267eded7852b34df5408569ac4191ee2d99b3ae30d88",
      x"0347bdde7445a04b8a7f001cc185b153be41b65f89092b4f0b7ce8574f20a241",
      x"2c77095b46de37a081d4299dd0d827afdad1d42db058d03d79cda6d5d3499b62",
      x"f04d7827976e5ff84ecf9d33bbbf3cc887af9b172216fd81b118ba4894de3f3a",
      x"5dc8b4df420feb7460e185e46a2942d3eed5fbf487efe657570ef80e45ab3b9b",
      x"54e356254db49eaa6d900cf5af286581f0c84feeaf29915ae0308f68a52f20fa",
      x"b4f001cd4a8d6729f87119807b904bc19fafcf6a9b22b9071efbf7d787631217",
      x"7266bbb5fa0f65acce11cf2629f13d025d585a2e6c0177780089f7ee02f55356",
      x"0da58928f3d020f629b77d8707d4bc746f46697d49d486c96249c3eaba85aa97",
      x"e72d46ac662df7b9c8c7aafc46b2d8da86d5d42052360d67d0e82eaa6503f47d",
      x"bc97877869a04505e384ae413201e8b2d2e128c6eeaee3b872d4929b594303ed",
      x"2ad5858a7e203397a9e092db644a0b1013025f7b5a3ef536c7b0d5c464ab5f40",
      x"0883a4ce17954cd7d06737740202b929a3ea1a9342292b226cc9a04b804b4ab5",
      x"88d6f4fdfe44b5e4ec55574fdf2a4a9fd4a5369d9bf825a3b40ed05f0188eaa3",
      x"9277658beab3da4a1df11ca0035b5297f748df236c6d4855eee3b94a2f17798b",
      x"370e38a036b4f86fed031a4b870d4db4a11c26dd6f5b89cd54711208ed02eaab",
      x"637d701e435b8d2ead8fb46a821efc85450e6d418543611252682bebc2c15bab",
      x"9cedf01be57b7b0938a52a0bc09741e8fab24049916a34dd9d1b93b53244777d",
      x"74d1cb3b92a7d0a7297ea2e7d9d0c5c7aeb0832803746f155b88c14a9d2c4426",
      x"58b789aa741fbf83eea74324e72af9acecd8ade8b550489ca8d8f6b49e10d2b8",
      x"69b63ecac50793eb7d7acc2368d1e240865e7e1ecab638d477bbccd7ba2f936e",
      x"401e23edc133084db1970aa86eb839ed258e387a6989beb631a8f11980a1996f",
      x"397939a8d96b54752e9466ac3a0e1f54537737f61a084cf637198af298f918b6",
      x"bc3efe208cc997438b0cda904b917ce99d0c3623945512ebc02d8346316e3c62",
      x"8be1fc19d3a54c53ad3235027b1c471d021648561524ae7ff027372c10ad78a2",
      x"8eca1adb707c5b2e7d1ecd6a7fcde96a43b2051769a7acb9f959455afa27b414",
      x"75eab7101e8f57b63770bc7c161e79f08f0bdc91b3386ab7b061c2185cd775e6",
      x"a898e717a4de7aff78d62067262fb68a960e3431d96dc131752ee6b95e9b14b0",
      x"b5ee6a3ac26b2d05367385b28c42e8d15edc5306d612c6267f87cfec8a0e9851",
      x"56c4ce6f45b4b18f8f7652d429a2b4f32adec5104794f7f8ca1179e74c212012",
      x"a626fea1cde20026c71bf533f569d0610603c5277372b45ef217f7bd7d5a6f59",
      x"76dd5fc45ca1b805bdf669cb57b821a0927b65d109dc2bf56b5358c53a589f7e",
      x"e14d6e44b313746f1330ded29489c1fc3b295e8ce2753571f7ebaf679cb428e9",
      x"65f0cad7c97af8618d9519a078101c625498feb3d0b139c992c420010a891dcd",
      x"85a785a960faea0b7a55a499a6c641ec63fba362e6a78a83e8cd85a7f8998fb3",
      x"5ee0e2930b7838289cd1c5a0f11c1f8c7d2a95a466c348f8d2aa1af2fb6f98ff",
      x"9c88df8dc956a742c0586d071228d384ec1e2336c2166820441f138f606f556b",
      x"a3ba30f2ce465966f7981f4628a1d526804d944aa949806a1c9269eb6da925e0",
      x"73e45f83f0725ba8bb30e9a2673de717062fc2f94ace65d4a4ae3295c5ea873f",
      x"12dd97a64a9852a2eea475c20d44171f8481dbdc8e0e4f449ec5be8975c4fbd7",
      x"cdb26fa36a70230804c1d52cc1acfc16b602f27f3389f91dd3da7f3c596430ba",
      x"b0623001271ade3955e00185f9cbe8c04392b3510de7b5a6a3a1b2a3c07f6bd6",
      x"fc735af1c297f53031ceee4417bf4665ab4945e552a08ae5dffb2c600dbd4bec",
      x"af8c548190b554051dffca34dd5c0555762ffb356c1ef86c49b3a535a7eb1847",
      x"c0d6e183e7a8018927b5c865012ce4a01693317ac2dbcb265aa096aa2e58d7b9",
      x"f85d8023696dd5e69f0c5dec1ff91c8ae57c49d2393d7a9e7bf6fac7f23f10c0",
      x"c8a9356482ee67a89f0a3b63b28b3b023b0914af21fa6dbf626f89a068747d9c",
      x"a30a2b1b51d415378648f5fe957c41720b13725fd568e78fecc01e9ef2165b9b",
      x"c8235f6b1773128cae03f728a50d2afee7b8e5468927129fb6e01870ca2b66e1",
      x"130d4a8823c0aeeb249ca951f98ab5a0fe334e11e2f078a806ddb492e73799cd",
      x"596d921e61972ef47b15a01158bd20fb65561bded50771837f79e45808ab2807",
      x"8e4ae6519e7e6237a934d9e3fc5613be1ddf4e84130fdba178e1adc3843e691e",
      x"03d20779f845f316de254888d612fa46b7b28c36ca82335beaa2d8af6d0c7137",
      x"086c696657d126705d3d14d822fe6b1a37d7de3770d1d1fc5d799854ff572aae",
      x"abe65de0ebdd6fce912a6d575f27fe09c0b0c350f10e45abd97980d7da3ddc3e",
      x"89efa6104f4a971e37c8182b54bdd62ac9b88affe088422d4698a2c9b15e078f",
      x"6ebbdd6f8e4e1c8bbf1378ec80dd87d29dc62eeebaa55e63fa3f019a30e386ef",
      x"6fb2c5be1dfbbd153be7bd26dfa5ecd3f8f74114bb3e77051a02eadddcd991f5",
      x"0630709124468d34657351e021becac15fbf3d252c911fa01f1cbcfb49aeb0a9",
      x"f53e08b77c11b5c1c90d44b878959c43dbb1f94bd0dd3bb159a79d036cd0b823",
      x"0c396db4a3fc252a15e10e0c0fe311246e724460452f258443052a7d51fd0311",
      x"6aca640e255cd4b7ca7ef6d9e8c377344fb7f8ad0ecd81e54113950f772e6051",
      x"2684ad108d269cbb780b698f61df3a3f3ae99197ad888050e7080bd3a2ef8d15",
      x"e55880b3b8dacb122dec9a4d2642f4ed4759508de541c109179d213f33d458c1",
      x"6ddcb8f376d13a5b59669fa1d372012837cbc1814cb70529f228dcd88b342706"
    ),
    (
      x"aed5093e61a7e4cd1c00c124abca3983a01b5789eb84bb3b54f4f594d00e7b88",
      x"91b72af920aafe3319ab72425d2bc09b1d53a0ccfb12304677b111c96e6e50f9",
      x"fb29a142ed0ab0e6211c823881efb479fb6565596a9e3a8deeb02cd82e08f549",
      x"cb00a791cc6d456d058fd9c9235e2b0fbebcda5c993a597c2c0937c21de04077",
      x"effcea1530f35ef973983f3fe589462c1dc4ffa95bca1e7881f0698c65180c88",
      x"c5fa942871ff4a28641a2c09d45969cc500c03b1d108a8cf4ae08884778ae5b6",
      x"a5b566e069557c533c89e6472d858a6664fda203ddf540f6149912828b609574",
      x"3358a109943e34056ace72988d40f19f6c1ea4eeaacd91c065763783aae8c3c9",
      x"26852df996d00a6da712383ffbb9dfcf04d08d52b51c56603f0c51cb67a61c6e",
      x"c6ed4074075b3e45b6b85e1e5dbc14534324ea04d21086212297e76674756dd5",
      x"170eb003ac505615a1452c50ca0f4e4cd07a3d7c4946f78a2bf4927971ce16ae",
      x"05e606234ccc43ed2ac326c8870ee715823f68f7c99a974717f2b589880fd347",
      x"1a1262d0d03035df3d55a80e3ebac656dcd8c756d2fa66e26e1da80a5fc9485d",
      x"85c8b8ea648784af2558e863d288a37a76ebfd00c3bbebf6332a0977211e5ea6",
      x"bdc7cafe101bc2018712e3deb72d6106b95301a34f4e6efa8e7ed0b85f365428",
      x"d432cfe697fe725624c988858821a621ebfd2c5929b0dc1b02f4e9358fa40ae2",
      x"ff34c4d4545f999426073c95e311f978f31180d4c65f0541a9c488f6304ae069",
      x"b11ea45436fd4f4e0cb7c1ee270b8817d7623ce4513ce572e94d421d311199df",
      x"2257e4d412b87db7e76a12af9df3e173813ca9e1a0a8320791c48584efdeec38",
      x"a0f3cb58c3cf5d51472f4bc9e04645c743852c572057d1c38219e5f5b562b902",
      x"7ee796eb500c9ce765997aa9ceeb7372303f10ce2e4598877c522023546d647c",
      x"96b7501692ea5f4f4a1905c77dcb93b16b25eea77ae7ec7e89e4eaf6c8a77fce",
      x"4faf711b9c3c219ef1f548ca426d523664b9dde41a7355719cb7ab8fcd1027dd",
      x"ddf6bbf412f9f1e1271eda81cfd1796e08266e7b8e8bcb59ffa4341d5218bf52",
      x"db81ab66d7fe134a21f7a85ef40eaa3deeb28a3372c5cd3d074c136adc2228b6",
      x"98392e28c0bc844c9618b6a9c4e665a8729082796ddebc1d93d8136946fee9bf",
      x"362d29acdb1d1a702dc3a19272284f7c404839c4593b3fa64e6e05602f55f9f8",
      x"21ecbd58eb0a5cb44198f07cad6e3cfdce7e8ff2844efca432dcbbd0a697659f",
      x"e597f37f506aa27713d22e2d5bbd3ac86ca03dd7c45555227258ff9929691b7b",
      x"2b16a425c3eab45c04cc8a0bb2285b17b69b792eac205fbdbad54e23b07d26a0",
      x"b6adf5094e0915cba6d14ed04a6f9215341de7613209f6bd7294c2dddaa4a51a",
      x"236652d3ddaebb202b51d1dfda5884bfb53251fceb206d2ec8728b78e5359369",
      x"85c8bd6178320e9e67004368b8da68c1eb917262ad33570e2060f523d3266794",
      x"422a2032d3b7b67d1c11dc155629d3a8d66da246021104fe3b97ff66cf68ee4c",
      x"8964c442e6820f545d2d0cf8f0b9cdfc2312913d70d586fb7b15134c20caf7b5",
      x"4552e9755f003edd368fb2cddc09277d9120f946e54508b344c1bdb9d5ecacdb",
      x"f940762b5e5ca021b7c2caec2c4325933fe1feb766cce5022f40b257c57ad786",
      x"2a4f79c17fe681197fb034998de633b404f9d2b44101cf8099ba76e555f8675a",
      x"e975a4e73d100a283d4d2ae3776d3c3622c387e52b1a93319361cd983aeebee0",
      x"ea30da5cd3104b4d1f5ea1fcb6e47de048ad1563605f89faaecadbe6b41863a3",
      x"01d2442980ed571972d142f20e0d3cefb87aa7923f92fb61077823d4a73fbf16",
      x"a5ead2808197e920b50cf1ed1cff7551fcadee5fcb9025703cee96bf142b2c52",
      x"69fe1ba1a887df5f8d80d8d5679d284efc4a0ba3c804bacadaafc53a96671016",
      x"5b2261d91a3f5eeb5b44f22b88db774beefefe4d639e77a8ad62b70761a59700",
      x"65c8b571bf328b2c9a676cba3aea403792b4394aaa066d5221c4a506be0fb460",
      x"ab6e0e42371a43b8887c4744159af082508e56590e9aae7a71e2c9fbb73f51fb",
      x"ddb174b96f2adf464a3489f9728f0dcaf9789cc84492ccf6b90e51a02f1e864a",
      x"59dce99880f5c7bb559cc5f62e9634399bc2bf7727689935a61a57fa7eaa1f8f",
      x"5a046ec9b19ca639b94ee7e3e7cd0015aceb63100562f444afd9baae1f18f20c",
      x"aeafe5ee219edda347ec8599c21725ad5e8bd59bf669e685bfedb12fbd6282d8",
      x"8723437835fe4461334f060011e65a6b2ddf566fc3ca4e4c706b90404e11b9a0",
      x"525d3783e1678924852270beb8a0cf9d2a141670e8682f7320574707a3e766be",
      x"07b7bc45ceaaf56bf151b9e8187d43d1b952db9e4e9bc626df67e561f6f5bd3f",
      x"10135abd923dc6487876cf17958b09c4e82531bf63efb6e9eb401c1e3dd654d2",
      x"edc25c4bf3290cbca289a15f45b04db683a4dac7dfcde6805a5d054122e8b2cc",
      x"dafb50cf8295f459d12268f9495407aced76d9d41b65c5f033178ce79518b4ff",
      x"217fcfe673bcbc24d238d0604a4cb16ffb2f0d580a043b47edf46439be91f4bf",
      x"e0722270d6bd47ea558f1ff0bdde7b5f6cfa377e1d16442f6fbaa3bb39cfcdf3",
      x"69a8ac4ec729b0d4d552335bfea4f1bc0b13cbf48a765b21881580370ebf6eeb",
      x"5c86b22fb6a6aaf2928fd5bdcac42a63be78655691f0f6e96b53229dc2f1bfca",
      x"25312b43e2e694a2bfb19f9793bb21d7e1c8f7a326cff38b9d2660b02460021c",
      x"f83dc4ebdcce2127f5b879ecf72e835441ae15e114237bb999faea60c6590fc3",
      x"719bd08bd17045a363e071b54fd813b161d8364789da97efa78ff4b3439c5403",
      x"507832468a85088fa290eace43cf8d016da878c154429e3a06a33e36d2e0b6e1",
      x"8c7ee2f4a00966071729fb2ffa9870d4ef74893718a84630babbf999e70952c7",
      x"b47115c7ff637007f11940c35b41e58611d94766d699302a960883a40ced1bdf",
      x"1716263b790a4128b44617299f6d6f0625b19892dcaab1540605b39a91987368",
      x"6aa353ae9a8f919694c000a07a5b03aa8935bced645bff1af3e51fb3922b0019",
      x"d7cb30f37c837c354c61f4737a9c983e52709aecee2a65e62a0f16afbfafe1ca",
      x"4f84dbc809e6d9eebbacf3d94984c39d2f7c2166f5f797ba63051c3454aaaf67",
      x"c702ff8876e0bc97967a22df8dc97a253a6154cf9fcf3816ff1a765905b7a019",
      x"fce29c664524d96b7d12657ab52172ec5a440ccbc2092a957430cdcd46167100",
      x"58d400f5b5e66c70e791942d60409ff9b94ff8b8ca72ff127cde4d2de7951f78",
      x"80f7ac6692e77d8656883240a81618eebb5294fb067a6279df0426dcdbb56049",
      x"03061a49d058d8ad98beb605614007caa6b549b10ac959480b3be6a7230d374e",
      x"5a0223a15d88624bd37c83bd6dd570757d0dd6390f1c15724a02c04b10b6ac2e",
      x"d28c648191dcd33066d10aeaf3a6f2ef16dca0e03c74cb2fb155ecea5febd6a0",
      x"9f7b66065bac8b13f54fc254d099d71086947c50e50560adb454fa2e8e129fea",
      x"14d6fad7cd6003c06df8051b50e9b902ba9df47828b1322b314c36567b9f0363",
      x"a6723555ed710fa3284102de6d88e443b0e878d0035688264abda2eb7328e092",
      x"8d6ea2f6dd28c5ba6ce4e99a8942ffcc20f86f175ec7700647a1f79d97aa310b",
      x"99138f4cdb4e8cfacce180f8f9507804c036a0fd52f8ffc86224297d2737f95f",
      x"4e42418f7514bc983e36fe6c0255c4e82acff83962110088b16d0f401df0f6d0",
      x"87477a61d826546d4aa940f6e913003fef405dcaaa7043b1af29eb25b88eb97b",
      x"68aa44ae46bbed6c3e6e69509a6a2902dc4e7731e90e1e5a270180698004c84f",
      x"e522c7ceee1943b36f1caea241cc36a66e4ddd19cd78a35681cfbdc290de10c7",
      x"3d04f46de1a905d05d672fd4ecd365ae3bce8f9e3d754fcbd4de6911100f264b",
      x"4c991eeb411d48b2d80856a1ef1422808e4b6e905fe1b1a7597b4f0e870bc7aa",
      x"d6c0c84491961a1b9ef81e25433c18ec4d9fa5e05d725e87bf9aaf818b8e727a",
      x"0e18134fac9f93d6bba7e8fa246fca4fdaaaecd18d9eb1bc38f1a499c5d036d9",
      x"4cdd0a81d4d08297e8aed5c527883c3cd8129e772d4fd8a40043e4728112f533",
      x"dc4b2695566a361572fad23f5eb2626cf1f179240d5d0ca54aa69661c5a93a8c",
      x"ee970e58123e43fa8677ba4bf448e7c3573574605c1e5e4eef357a6c71efaf7e",
      x"4fb42aabd7a5779f82c6936ed35a773bae8d72d209f83aef5981cfbdc65a5fde",
      x"fadd41b8cd225fab7b593bbdbd636006b27cafbccd9bc9a25e4a19481fbd8282",
      x"92c609632148c166f1ec0b6c1c1cc597e1f73a9590b2f34c2c6b9ab1cb17b576",
      x"c94e71bfc0e5aba3fae27051670fa050db2d59245cbf5739831ac9ba44838feb",
      x"bbd7f8c194f1fe7af09937114e7944d9a6f268b46fcb24c9ef2d9c23e4f2c1b4",
      x"a28cf0692e21bd17bd21da7325bae0bae71d10cbedeac9877a288347ba3a5a4e",
      x"939493bb2f052a23380770df0fcc69be66f8da6ddd1c65836597a8884dffbfad",
      x"e1459025333d9463068560a6caaf486093ad1f83deaefca2b3677bb5fdfd61ac",
      x"a480738cd58018a484059854f14a9ebe733bbd65cfa739172cb39bddfdd2ce4e",
      x"2d0b6f12343940466e4c7e6531b0318451370bed80acf11ff963bd7e90ceaa16",
      x"d29f0c503edc860609ea82656e38f90c5c189b4061e619ff6986e175c43fc795",
      x"34a91d13c1111456fbe8bdc601eb60cf39e6a9236a1ff5a54415ca895811a38e",
      x"3f83ab54012773f5cb14534decd2f964026488a6ddeca2f312f79e3cc5ab7323",
      x"02d8e980e972adfbc36c5224c27d388314d74ab85fc9cf00688e67c94fe194c5",
      x"accbe4e2b53de068f91e89376b6af26528cc79a6df0990b3b37da91c61186bf9",
      x"2b82922163b26c53be3fef692fbf00925154101d1153199da278de3f49be0d33",
      x"d9be427ce4d17de870c4da60ccc2470062694f87cfa2b8788c4b3d66bde6249c",
      x"d68fb852fa834dea484142b96d26878a5cb2dca2da78734b7068086c7d94fb85",
      x"ebce7481d119273a4ab47e6f23dd1b9442054a25d48400819c1513a5bd282ea3",
      x"b15e617487fc9bb3d9a1b835eb5ce1530bd4b915f72d9f2d49c84ce32ca31670",
      x"408f6c1757ab9ee58c0c203998ab032bd2c5aeb03f527b83ebac0f1c0af7eb10",
      x"1ab4d22182832c915656f216f47e0165eb3c6ffe74733befbf1218e07796448f",
      x"2b19fb083c57f124b78c9de773de242615637c2186135c7e119add005052565c",
      x"9bf49ed07b66f88fce8133f6b8dbaf722939a624486387eac7edff1011e25b08",
      x"c0778c5719c7fbdf7104c18e093c22b7687d7315abf62869060baa82f0698f50",
      x"72bfe7b2ce608a748b5d6519828f6a1bb30761a11c3610172545bae7d1412d91",
      x"f7f14ef3d2cdeaf26bcaa5a0be574a45db549fda5e576f217083f749c986492b",
      x"aa25aaf599f4c7bc689612fe7b148ef9d8c4e45b9cd2b23a348bef920824f702",
      x"5ec58ca5b7caeb176693afaf983634aa766ffa40425833471cf4a5498b99b2e7",
      x"c09c2c3e85bb57eb4aeb6338c83cefdf33fcad1592b769c9f7c0a8773c6603c7",
      x"af8e409209a348b393c0d5c77cfc55b8efe9d07a9c88b91d38b7a6bf719e780d",
      x"5cba0fb8daaab38c56a07a918374433f9f43d7a521621e7624374f86b23c432a",
      x"b10aa975b5ce35e2b7da8fd85f312905dee947325f437959d54cb011a467770c",
      x"3cccaa3be5f63957ea17634e1be319b4c39a289d276a26c4dd55c01703915470",
      x"b52f9a257d75939e992dc99faefe04c2c5d487a8705aa9a7d75cddbca5867210",
      x"fd184d6a23f5740aa802b76929d4a2455639a6df536ab6d3adfdaa8f131d4ab0",
      x"0832376f3d08bf3bdc4802c5661ba8f666da694640005aa7d64c5af60c71675d",
      x"8f109fb5022717f695314a3312b3f2ee5a485290d3ca2db0f68cbd0c7547c671",
      x"bf74ef7d969cadb7da068bc53e781bfaa28a378334e753bc64671149be5eb155",
      x"18b5629abce0f54a164abd51febe3ea6599185606bebf08e8aec3f526a19847d",
      x"35238244df65e6b78751576f9e1bfd419f76ea66cb62e2cb4c07228474de3058",
      x"cfc69026125a6660287c332aed495adf2c0e0c62bc409349f923273116c6ce85",
      x"ab588e8b90a8b87bba14b3947f979f98216f1551afd383dfb78646fe7a07d2fe",
      x"e5b21304688050ae6cc4534cd6c539042b5b959613c8d980f7dd608b06df433d",
      x"60f9d42c76c4bb9a10cb6c0a89526fea235f4bbf64b2f5feaa4f3c4b03e9db7b",
      x"249204c3144aa2f6217bf846a945268a67bf5873f1c82f35ebe28a3e350d27ba",
      x"c7a2633772491d514837763868118560ce3e9b008b1f906a92ec280567bc707c",
      x"60b6b2623a856b83faaabf2b48d60df875bbac4b86e3590b6247aeecea08856c",
      x"bc2a5317856b33f5662a55e78892d1b3a688080a4ea159671c39a211da0d5874",
      x"b72a40042707309c3892e25fc2b8080d500fa61940082aef363ed0ad03d7651f",
      x"f8d5f0bc1b031bd1bfd3c729779ad6098b45edc4c341dd92fc74ec6e76637752",
      x"ed4ae5b512650f8825c38006a0530068bd2739e442446de0bcb9a2c2bc3de866",
      x"c90494db399e5362ae3ad13ed5fada9abe847ded428ec2634c7d608f363e3b4b",
      x"2375d5e678d6826629962b1c2b336164c695a31f0220234d7a2fd4bb837689a1",
      x"a37419c7c9ab760751ef67f73db6ae1aa398d6e0d6fd240910e4f357d92aeb4b",
      x"c4960e8730b7985737b40e495cf69e54409d2cea153f8d6a9298736ea2339b13",
      x"27447ec6a936d5bf7347f3298477d9129a2424596eb716b44eb86e12bc790bf4",
      x"9ba58d81c19d1cc536968259d9e4d2e2ee998937b8d2f45cb14c1265b25f0a06",
      x"67ee1c4d384471e68537b750b72dca7d22e7275b78503b3fc136f45dc8c458e6",
      x"2e4d34fe0f8a03f982d630449463d7e2ce7b32cf9ac86e4dae95cfc7727281b5",
      x"74d80bbbb350c33572f0168912ae67933d7b30a98ebaf27c168b47f2fc69c4da",
      x"f245ec7efc55052cdcb01fbca66bc0d6df85a9e2ca70d1012cedc9cb1dd2495e",
      x"d51f0a38100601723b101602aa96a7db54ecc26d9a73c401fbbd755d480f46b3",
      x"70e88ea276ceffeb10a96c6ed420141b81f2b0e6cefa6a06c03c5ef73308091b",
      x"3febdf4e32e017b43054afe5fa19fd2c2af3e137e194c38c37e9812967737f66",
      x"a1e0ecffc4648d069d3b104c3799d4fdc33ca85c8806f775922eb4fe58fca003",
      x"a0fe5995c7083af86945e9c46216c727173b0806141abd39e9e0b778b51d0357",
      x"e34ec1f7abdf7547bc83374daac500a9825425b1ffe4e44a44e9fbd6926b8f40",
      x"1df36c4e1bd639964615ccfc331bf3ce2c628b05404bf69fb1ba3e195d556aa9",
      x"734646d8beb47db223169ab22a80da9388bc5cec1e8f00abefb38e8f4e800f2e",
      x"3771a7615a85d3b790ab2c533cb4c17ee7723a30041f728057d2cd0460efc052",
      x"873ae0dac3b60b65457c4ad6d53be5c2060a03b78e19c51c1347e50b6ce59001",
      x"17598dfdd83e7355f883511544d98d7d756d692e8e8386e358a3631259d80abf",
      x"1738ea985a061de2477b1806db35cfb5e25f2d1b4f601e05c954384a5fb33150",
      x"5c053c26a8cbebe54ef933d87dd31302d76d2e46bfdcb7fc6f1c550f27e37952",
      x"40bd143b29754a4623bfe67ca2133e2bd03a7b1842865359730a73884ccca563",
      x"4ba41faad0012e372075e7451686b1de89e4e8ec6c1a6f7b1f5fe1c15fe02202",
      x"b0d0d286b4d0aa17001de69ca7ef9b57dd47caf3de593ac017163622c6f24976",
      x"4b605eb60ec0e9a1b532eeba8cc97b97ec923621bfe643cd75c52119ed60eb51",
      x"30aa8c426f11863a07966de0cd586857190be5a25fe1ec82d3bb1d8efcab99f0",
      x"4d8e8f53703c51b534ade556634642d6f131851afaae15ef393fb54b0ad6f3e5",
      x"05b9c8be48f974aa79caeba338586c09c7d1a2b66edd49f016c70cd7933dcabf",
      x"f81a4396a9046d5c0092fd29ebeca7350ed97bb8f87203c4f67f825a203829b5",
      x"7e2d1d2a8265863d8a87c2315c92edecf5a99d29d78d2a39a11522d54d9ad57b",
      x"39a0ffc674b1046da0cc588212025c4c777fd2253f75455ce10fee1ef5bd9afa",
      x"17fb5fd9ea989523470d32da0a53cd23ff49998c5d8d76eb000f1a11b3306c0b",
      x"fd963a4e6de8936cfa0811640286462207f2e0e7247756a0539cbccb6a7ed4d5",
      x"6f20fe6917d9eda190916b29ffd5ac8909f4b766f383b766a2206c747bc2e36e",
      x"ed20846ca0706ddb42241590ccc7f81b877394a60f897d7e6fa496550faef251",
      x"853686d2292d37ae45c90e5b77f4dfe4a26b8cb728c31a3f107d2b7be5d46c6b",
      x"7265943167c36a9f53de42d59ff5ef1bd21de4687cad1732eb6ff6e13e420a12",
      x"108a626e205e953ed0ffb45ae8e55ea4e2d6f08007d84700b42e82ce800fe1b4",
      x"8e0499aea9126e5f4ca1803fc4d67ffe7055a692fb311c0dd19637475f2f848a",
      x"8628d173b8a9c45bde5b829c29bacb5e1707786b372a9e2615e3e198dbbb08fb",
      x"5545e089df36668126e68eed99ad4b347e5726f4b8a1b13ed85b4f6f17f85c72",
      x"921070f740461cfcd6e80b163ba1fedba0a457c89fd5f5e53249eccced3438db",
      x"f5046749973b1e2d1b4c3f4c15dee4189aa23913c0b5de3e9d806fdba16a6371",
      x"c3c5c7464890fcf71cac5587ed5907d486de8ff6af626ea12d92ede504df1c35",
      x"e7bec33148a63b45194b719a15897c13d65db5639cb78ef987f64e3e014e8765",
      x"fef31f568ac1f89446e5a2e2d8247c8545384576f7c8287742e459c1fb97642f",
      x"136c68a149ba7bc7e9d940702a0a913504e5339bee95b4f71d6b04716a2721f5",
      x"65c95b6b249c0b9c8cfbbef33709fe424ac28327090627e3e589b0daee1695fa",
      x"394792c2cef193f92b0c5964e94147b41d6ea9a5692bcd2bda6cf1ebe8617763",
      x"18ccca75d71fce3b4e005ce7d0c684166c89dcd1857240aa7e1022f0601ea36f",
      x"4137b467b6ce5f44b639163860669706408c8cbb1d517ec920fda0e3061f6fd9",
      x"bf8a5a21fa63b64f3c9b66256649271f58e6d87cfd136dfc854a35895e028730",
      x"62ec67e0a417d463851a3e8be6a496335f80bd8fd62c5325349e358bbe92a4d4",
      x"1006fda7086174528dce569960453a3755a1ecef294db6e90402185eafdabc46",
      x"97e23efebc0565b8a869b37ed973f6b787717cb0b15b0b3d279f8d000d5ccac3",
      x"0dd05178aa6a4d892359b55ef151fd831b5ef4b2101d2532c0da123b431c1fef",
      x"45993f3b50714578a1e68b44df3af2c19146698ec7fb7f6d37c0b41254498928",
      x"59261052cc3df2946b9f749fad9da966830ec0f2d78e4ff99aa11716be4c5b83",
      x"de62db719ab4b6d8a9c29f4757860504d856dc0d2dedfd698dd274e9bd95517e",
      x"a0dae4547ee3175343da46466d544a22bd637e3a662dec36cb653cda3b5eea8d",
      x"19586f038c23dd9ea74f0b06ccea2d233a5348f11964c83e64752777f4390890",
      x"6925e436aea69fa58fc836aea8356a4c9039d8883c1c7206ed979b2b9a5bb7d8",
      x"9ed0278231d9a00abeccede1761436893c58214effad6d8b6b70b173835e0e53",
      x"9a6de3e6ae1e469f0d7c93afcfb8e166aa1f59aee5dabcfd5dc9c627d42c0486",
      x"567af934b2133984efc1373cb79a46bff5a953e35adcca46160d42b17b3c2a2b",
      x"425935bd7fed747f32aa4b7ada835d9b21209602b9b762daa55dbd4f2152086f",
      x"ba6d625959c5d71e24b8440a26003c0ac255b3c63df7e7b24192582697f3f922",
      x"9c7ff8c5a55b195eebf51d162d5fa682e419f3f2cd4d454457d177807d6eae88",
      x"b68356d4f6b2635b766dbb99ef5fb724bdb80d3189ce779fcf3d7588009c48ae",
      x"71164bd236d0a6638595cc41f99967b9284fef4881e65d8a8658c04cdd78f129",
      x"fdb3b984a81fb97ba943af45a27e52fd396a2f6246b3662d486ed0c5de0b8e7a",
      x"a65bcf3d97282eaf19228a007fd23a4162846cf34cbf677a74bf1288cad67d99",
      x"504a980cf0c7a91d7df6513101684d83767379feabff651e9526e8dc04da8cad",
      x"11ff4f98c5a638810d95fb4d3fa79a59d24dfe828f15467fcbc440deab638e5c",
      x"4261f8d834f3010451b4d470902702edfb81076a6c99d87ca145d9d43f3f99e2",
      x"4c749a851ed8a794d8742edfbeb6b75f3bc65904d54f18e846c76d32ca0c3f9a",
      x"8f278e34e2a392906c51fc68045582ac32aa73b5607c58180bea37ed2b16def0",
      x"e833360e2c5c627e7ce509b962782ba7c82fded0e5cea98052ba63afac3f7870",
      x"7c56a83fe943c97a7d6d092203812301b670dd86a0414be4fa2c57cd2ba88589",
      x"1815333b6b341a0631d53fa11966f8428e3a1b85b05114c7dfe4c7e6ba0846e6",
      x"035f429132aa6d8ddd8f22eeca228a3d2888f850f91315d83fb762b5c6314915",
      x"390281b53921d175d519ce91003e603783f9ffd7a0af3fa78e00769b65dade57",
      x"e22afb560316d4000fc50744c54731d82d8559219616fe4bf567048e7ad04b11",
      x"e16054452053d05d3ba20b181f47c51992b61d1607ccd28d5a752598a0d15bf6",
      x"8376a952fa46afff0eeb600170355cf903cef89085b4ef711ba36dea0630285b",
      x"20f4cbb58ebba98022c3e3dc47993997b7b71df107a9c2937a7be1d03047bf0b",
      x"8bd192d49a9fde7a76b27c1cf22e7e6c055a2cf1003360fce77a60f6092b09ba",
      x"a2853c664e3153307e899da03c1b8ae45adb106693828c33134f671132f6579f",
      x"ee4ea6975a9eaa318e2fae513306ca913bb49336c2fb2c6e6dedc30083e52c00",
      x"d6eed5d90f247ec1a7ef7c0d704cb6d047f236715c5dbe72a5ab6129f79cccfa",
      x"59acdc0fc574e96720f808e781057ffa6f1bc7447ec7b18562f1d7e624accfba",
      x"eba55f55ea11e152a7870d34abab319a83089229fa37c8573d9ba780564fe5af",
      x"d7dfaf3a880cbde6cddf331c6e0f7d09cecb60cb456fe77d0323ffe9b05b67f4",
      x"10459758c11ae4849d619bede075362fb799a351be30f819f786003395f8c6e5",
      x"c925637529736b1f520607ed73860f9de57868a81ca45d60d9abf142dfe01b2e",
      x"9442fde0a1d42614a55ad2a6dd2362c2f6db108ea53663362b42faed50176c0e",
      x"a797dc31d0657de1fad0e9bed3db7ae02a9940c79ffe32a6aa4c6d60a9fa8db8",
      x"40aa4ccd7ff48582901b3053a356ee13b5c51493011ffa691640e20ea18dcf02",
      x"2317d2baaacd086a72d77cb1f81f327893726b123cf09dadb1c07b2b2956b138",
      x"14f72a5c66c81e7b07fa92c8f451a92e99aeb29605ca8b084607a428c08ce657",
      x"38aa769e34b2aa11381f037048131cc3b4983ddf65ac129256bba0118a7e8dcd",
      x"be44f5f9b81879d5c333571e7988b510d4e102b60495a28d16515998df284028",
      x"5d0a069fae5127a15e58b761f83419fa1011a19f789685084f7f1459426c338f",
      x"14e95ac3e2375e22ff3819bbcc7926ea289fe961dee3050429a3782c031c443a",
      x"3b43b9393665166d968bb1061aca030d332b95067161b98363914c6d6fc89cf0",
      x"e25e008033c3007cfc6c96a6dd27805f026c56671c6d7b73d898d92a5cb3151f",
      x"6d054e693e5da8586ae400c765233fff92d9f23a92a49f9b877d099f7043f358",
      x"58d16dbaa33bc450ec44ec514126eefe20952f31e1b2f2f64ff7ec56e86d0821",
      x"29baca6f5fc382e278286235040ee284cf3458f22b7a5d5c32430112395b7e6f"
    ),
    (
      x"6b4af557233f0112821398f10781fec3e1a8ff9406090f67bbbb61185550d11e",
      x"fa205c054d9abf7d82ffbeca383a47a4ef274c632858c2eeca6011796341bced",
      x"3f0a1b512ed0a4246faef321dbc14cb99bcb92b700bbc366579443cfa3789dee",
      x"883874c826cff422abc44fcaeef2170486daecc4dab6eeddf0dd104a33296225",
      x"db18c761bb938f5671794c32ffe859083af03df64ebdce25c93d5635c74a041c",
      x"08a88e64032dc6150cb8b16531d39e3771e1d6500125640fae395b8cd69b32e4",
      x"77ecd0cf647303f5d41d0d43adede7072c865a677046be01c5a8f59583719d00",
      x"9aa214d7ff3da2ef37bf9295ef870bde7cfb9cb3dbc1631fcf127e31f53d9039",
      x"9061cd85a3e5944924f9e6e91db3b7048af45cff7820d62a9e8b3137199c765c",
      x"2a014636cd10465e66c2bfd4f8adee59fee909d7cbe852ae46659d69e6169409",
      x"4f611fd65f4e7c6d5e3a5110cf1929ff0455d7b88dc509c2500270cf24945dc5",
      x"41c018f38166dcbf2f8cd2b047b379c34968dafc38d1e4c7f0454a4f93b77db3",
      x"8518ecb074434e79dc4803c52b145c204f1645d0c8b1f50d24804bd2560bf9e2",
      x"e5a6c70b786e3ae0f74fb8a1ab740eedbe53772b8276dc3298c7056a0fdd85f0",
      x"effb7b6852bfabd767c834af2e05826cb67c8c54c49d17c4cf8384a49df0835c",
      x"37f32b662025ae3682e64660988daecd6a7436cdadae2264f1309cb82e9ae27c",
      x"49194e082738823c681f8939837893e0e91bbaf824097f3f749f9c03b92e4749",
      x"06cb55f4c95421c1117aed879aa6815b13ae834b8631e6c8710d81cea75cb264",
      x"4df2b78c04530a1b87ac09a03971ed185c3021af1c260f48e78fd7d7e79bf789",
      x"b3a86fb13b5719f9d84b7dd4ed3cdeb6cbca85e3bc6b2c380083cd76e955f662",
      x"70a0d1070670a6e0401ab2ea64a9adf75cb659b1a3774563530614355ef86502",
      x"f49205cd524bea30c13205c7f3ec19020d3b040f7efd24fa82daec9f245e9d2e",
      x"58beeaca293017c0d3c3d92f8d60855ec82f83e23f1ccb10bb350f0d314921e9",
      x"1c05c8ca431480cdb11567598e3c499ea59eb294bc7cce122a88f1c0212509ee",
      x"dddffd6304735609e534a7168817aed2734d709f980159b0107c94fd80cc4f76",
      x"d6e31b20883e38a4e26c888d856d8d1b1c8544db5846445c40308bd3240bd896",
      x"892526a89934b5eb16f18227517ab18429e2a588bf0d261b46e75163f6c8e02d",
      x"aadd5e867dc28e81a6b93dca20788739a8f4bc7b19466a1e3439f80c3eba21dd",
      x"c3e4e0a2aa1af9c6e63bce833169091eb18f7efe0329c9ac97aeff8bf27caa5e",
      x"200920fd86071d5c972f6b28d3913d2c13f851d9beab4eb2a71fb72774d7ee32",
      x"8d296535765fb6f57f10db89679254e5ee3c20db915fc6d2cfa7ce18c2db5994",
      x"4217945c67aa4fff899000edd870b1f61bba64ea03886398094c0db675046371",
      x"a01bb4a9bcd88efc89ae6d761842823c25d761645e8e6f5d26aeb6812e2e7d24",
      x"6648d0575a962eb85961bcd592e7517948c713c27e45ff3fad20fd8c266f8ef7",
      x"03a76d998de9b8f77558e0fdfd80e3bae93e300a3da4a04a7b06f905c9e00194",
      x"ae55d05938b352b0e87a095be05fb48c5d756894ba3ca01d78810e221fd08874",
      x"01d7e9951dc89ae65ed8e459e3b9340d64a2d8ab91ef1c9b1f849e03f06c3557",
      x"8bfe7df079ac337f3c9ab788783f69732c64fe7789e64ee231d2989e5918ae03",
      x"11727b81a2c1b91716948b36c64027f814c424589e9bcb751173aa2d96fd24df",
      x"8604aaf996c926c52a9d10293342bd2849ee8b315743e90d3614a83c8f28c173",
      x"b08d26cfdc3afacc48f0e2bd7364f7b561f0170ec76069dd9a4f69a71c4cbb86",
      x"3853267aad1ec74d98744a3f04f5fbcfc7e043773b5ecd5b754da72ef3f74c9f",
      x"b92c6312cb75a0bdaf1f25c3b51b47a0d61d9472b8f520baaf4e7c6e9ed1d82c",
      x"99bbbe4d177b125c6ce42ca1625d189794a7d1491f7ff060689c9c3abba22442",
      x"5eef2bfd90bf105a24e87ddc6bbd9e400dc62610be4a0a46674788de901f28ef",
      x"9e79dc2f830b943b9ff31b61759ba355d50dbfbf00082d2311759cbad8c17a95",
      x"9c296168c8966eebbbceffd456a992b64f7d08a6407fc6e50e61a8546debe270",
      x"b0ecbee25b2454bab36454004463482c45916d8233f1fa09fc2f219117d16782",
      x"7e39c4b92748a4bef0d69bbb14a9fa832b20d6a661243c0034d69ff745291a4a",
      x"59ee11d5476f135c2db12b5a5bbd7e72d7305ab371c18a42f6cdbbe58d8be763",
      x"1b0fc75e16b9ffaeab61586e193c1faff5302f893e685aac3783b966fc55fd44",
      x"39d2a3fe086dd07c1691e0b56d994e5fddd68490e405a5970a280dc9a02c0c25",
      x"c7cf8df509cfba1cd3ab3935cf7fe1baf41f5503d4d18ba0abcc577f5fe745a9",
      x"9aa8f8a529599a90e0796ca6a13a0f4805901445acde51e310691941d51c22e8",
      x"d9c3d4d4f1f8dec58a364270757ad65bc0e704eb1d2ed675fb94d43f39b1d420",
      x"083afc7d00b78f13d5ba80fe787bebd44ad093d18c6dd440337afa02ece2956a",
      x"5924f83dc418d1580055ca11fd73a15820a5412234c36839df9c0ec38704af81",
      x"f5da7ca6f51273607e808c507078f5fc3a316085f8841728e30551e189200868",
      x"54703ab3a3d214f9b7734e753fa60bc853e5956de1d308208c91865c83694ba4",
      x"67071c7a20990278210765deef663abb38fdf434b09771f6fd32d990af13bada",
      x"271b328dae2f54f95b91778710e4234cdd48079d758ab166b812442685420d8a",
      x"77975a4e62ae057467d499f24c9a2ebcbb40131ef9b81e6a3dd30b246502d806",
      x"da1022f8f21dc2c269e16606c07ec81db746f19b568405b4198d0e928fc84aab",
      x"657851f2653046822b550dc46f509a59535f4f69c35700adf9c30458631d81dd",
      x"db7a0676ebd961ea85d8f62b532a4b43dffadc3aa0f4416bcdee09b3ba7d19cc",
      x"f7fc616bbc0242fa52bad332904c57d722c02403916fa45521547e6ecf54cf9b",
      x"a755bba0254d0946e2acd3e952de58c169d6b53c4b12d376e54fbb206afdd4b3",
      x"9a32067ef2f8ac1e69bd97efe8b8699736eef5f3a77526733c38c246bc4743d7",
      x"07a53ce80e21ba61de478a87f6cc888b14050f16c272361371fa813e4841b795",
      x"ce0597516ef9b0391333e1e6bf6285e7c159098153438ca635e4953f9ec7a20b",
      x"034c4220b6c17bca6a6d39eaf73f9c7a9d96fd867ce5c1347cb120205c123525",
      x"f8cec6298e3d86e4bd5e5fcd6c9ed20c4481ea4cbaa3f988fa96bd32caf8c585",
      x"58ed10d2b383ae4dde9989bf1e90ec9b03daf34004dd4252c81b0da2e16a1d09",
      x"37cfe9fd7d9a4765c2c2f4f44466f42975e487646e0372749842e910c24d64a1",
      x"fdbdf9a886db861e6976ada7aed1d494125e2628407c2554d6f963847fc94fe3",
      x"b1456716c76b6ad2e59320c1b099372640a6dd578d98e4ca4af83ebc75bdea6f",
      x"8bdc20e57f4c2f8b7df84f37c306cd59512fdfacb1abb01a9216544c8e9736af",
      x"06ae90b6e785e67ce2899bc5d11cb954f52ec1fc461cef877945e58233bd78f1",
      x"40dad6065ca4bdfd765068e2e750afbc922f75b98df16a51aab869fdad2f572a",
      x"3f5f85ea6e86d0e3aa5f95710b4c9a05dcafe1046433e2365a7b132b9ea30106",
      x"e5019a1298abac7a4f5242d8aeb8c1486abfedf4987ea0ff6062c026b815b0ca",
      x"614d0407df140af55dbba456b186c40b8ccf4b90c2ad03954a141bb67eb25ee3",
      x"2f5a84c5988c5ed8207b203160b9f5fb01a0e59e16f11f156a0c061c1d5502a3",
      x"39e187b460e708bf476f72245a3722a2233380fee1e0117d566873e8de3a4603",
      x"0cb86eefe714b7a57abb3bf16aeb70e87ac4325323fdb5b4d630ebf2a257a971",
      x"3d5752e4c42240205e4bf1cee19b3b04c2c694465451d9fc74c45f7614ca560f",
      x"94a1e5b58e27b00dd9572b482c9e9614f7d7fa6a3b4325261ba0bb3b54dd51e7",
      x"e7e5a90c34bb26cbfa5832009e48e6d296caced76a7ce10b2d162eadd5402752",
      x"729dbc62d62109439555d66cabffda6c5adeac8f33918a2e7bd91ebbbe3a1918",
      x"9c625a2f4fca84c86a2e2aaa093e8a71329cff78a5c973a42a7ade84d9a507c4",
      x"7a5dd387228200a1ca9c252ea7447e32b2557dd31588361acac3691de4e678bf",
      x"7a96a6b25585de3615dcfbf0e1729a444044bf42939107f915e065bb825674d8",
      x"07f1085453cbf27590c84b0ac62d8279835a2ccd4877a98e248f3728d62f4216",
      x"3fc62ff6e5a3c00becbb1af7fb4da4fc91cfea2c67fe4ae9e8a04f0d332c0d08",
      x"85afc505301a00228ffab7f3916c5eed9a3403806616a7c50f723b0587e36683",
      x"bd72b425920f52ac04482845e48d69c3c56988aed3070572bb94535f3036c5a4",
      x"c0408cf7aff20d0a037edcbf664bd17eabd241957f0489617d986943ea2853b7",
      x"f5e03c9b58604540fe9beb5291ade2ccf695845290069f25dd31b8b269578398",
      x"d16d8f0c87ef8e8ba911403f389cec18066a6e4451f97c536e8ec39ca690cd73",
      x"ab1a1353d3e7916f5225075de2bf97c7c9eaffa4630042853813effb4f6266d9",
      x"be60711384c41a96fe84a03f0a29779f6ce6266178ea8d3cc79428bc9afe5a35",
      x"d90f3f481fe88068ea26e97e0d384f82096197125a55e7388b0b21c1cfa4e881",
      x"67b6e6b0e43c8c2ba2575c6fb9375007b7c5c48eaf5e8936b749100ee8ef5c95",
      x"e4c168adc456d283bcddd87e5b25f6e706795ebf94d9cf7a1f2d1b513e559090",
      x"d92f229960efdfde090a4b937480b34bca431f68fb3d6a9f1531b39febe11d36",
      x"d9a784d3c9bfd713b87b1ab272b6eec9d6f27985e27f08d97ac5c432166fc17d",
      x"3b382414e1b5227ee7ba0a723e627fb41242788f17c764aafc8e9479cce32949",
      x"ab54262fee250ddd6741575108f56d394bd59696e8842d15b21d212abe8b1fb1",
      x"271b3229850aad16364a6fc602038894860da555609ff0e4f60572a643a8686d",
      x"01bbeaf32154c05f84f8825724b4d8bff9b876bbca78947de9ec2fff1f671a42",
      x"a0e6f612f936f1f130144908048cb554daadcc51272a1ff8fe4470817f962046",
      x"a6d1604887c7a968dbbb204777648ff977d1c9ee60f2955dd5b106394df34052",
      x"b9615d39c5b4befea7b4a919333cf56b2d43de35b77567e3fdec0e389628fe57",
      x"c548552f01d6c937cc8b31dfc17277cbfdd7e2f81581b6a16319e9a1f23911f8",
      x"6b3bb0c8d58690cd5e6912d4587bd82e29288abf0d8a61a264459b564f738aab",
      x"5234f46ef4fa6856e8c72b098bf1b306f779a7d5ecfca6ae1f1ec81c00ac138a",
      x"cad16d0d5a6c51ea4d89ae3b6be2dee09d2978eb96ea278f404e96a9c20e5130",
      x"d1b1b392f177aaded619bf382018ec36d60c74a20d611fb0ca948f32f20cc9f1",
      x"ee3dd34079c7862e49249aa376bcf88de216053941580ef8e084f0563eef8a0f",
      x"d63a6ea11b9959d428c77f54610fa8a049d84a62922a1a4186524ed2d9b68b56",
      x"a32b01d4f66fecbeadbab047225b052a8ae20985003eca0e5265a7aa3dfc38c6",
      x"074eb442d3c9bff8cff7201c9a949e6024dc053060563fe31cd17551820cd71e",
      x"a77f39911ed29a2ce375335167b807cd88c7ac09c40458140a3157b57888498b",
      x"e5fc18fdbdb2ecfffc0cfaf9e496ca6a3d7db5c64bee2414123a2b010deeca20",
      x"3a6b80e287b190fb8a4b13f2518ef7ff4dc4a5d5f64e05b1c36c739164e64dcb",
      x"ca8f1e6d6493885c587b9b8da43138ad38bf9447873644819d8a9a1ad5f10045",
      x"5fffbfc45147879e4146c48fdce30c1355f073e7169617f4c03a242ddc774703",
      x"80513205fd13fe516646ed9d259b34f510c224422293675acd0f02191fd14ea1",
      x"0eda4857923ac56ea9e3f55aec17a85a1e64a3b5c6ab6ec5ec215be3e961aade",
      x"a5daeb4f6c15fead26e6942c8d7c0a64243e3ee779a75692c882da63d1a51f51",
      x"e3d1ea09cbc123508972a01512b0dcb6546771951ecd5325537a74848b98c4eb",
      x"2cd3b836d3526d4daa0adc7e5cc32ab964ce310d7c061cb477984ca1ab6bbb8b",
      x"d7d234be44786f040a817b91ff3110ecf09f156af1a3e26169ff0f3dd97450de",
      x"449c882fc1da0bd77dc8982d52630b62cb75fdde3463b70a1a9f64494a41fc1a",
      x"e58974b4e15acd683c52fa0def22f8978f24bce71cd19ffa8988e0bd546ae14c",
      x"fe6464041ca804952b096f1e0c371f56c3ab980c6c55b4f5b65f3b64b56f5efc",
      x"1c22a7aa3487e1083a29bc77d54ce6deafd4bbed19e3aad6d768adfdf446e260",
      x"a3367674d0cbd9279007da9133eb60a2510a5f44c19db52b30d35cefd957979f",
      x"09c65a72a6681854f92bcbb2e12bff37589671e2286f6d7bcff2b7ff42d09353",
      x"e3c8f5075f656603b02831a0d6ac505fd011d1faf320c20a9debc7e7fcc18c39",
      x"eb3c8948c8cac075413346c94e15b12a889d04caee68cede676b2f3874d64312",
      x"5e002bdd731a6c10cb68608015f5b446f6411273fe520ec53b28c9b5cadb8d8b",
      x"1f3ad74f3399bdb46dea1bda8ef33812f8e7b9df3f86f286925148046daf5e6e",
      x"409f09e14bce6b4d1ba622c92a3a4fb696a155293999de45b407c6d992c75b01",
      x"7f77fe978564f0777a375d33d6a0ee7ff42116bff5d7c3eeb6304b76e87f9124",
      x"a9b6895a16c986d97f5abc51ac775b83c72b68db04fc35f866c346c47b3a851f",
      x"62a8df1320dc8fa3aae11926a591aaa0b1146bb32a787640a015e7a2e12734f1",
      x"b0658a8746b85c048ca6e6fa06db43b60c37eda08de2a4a4ad228ea81db4d366",
      x"a353c521d0287e8202a622f319b4e1820d2d1a54d128480d58696b8e45f170dc",
      x"d66f2a788576b499820e079b0551f9f8e68a1f87f8eb27d1ed3ac514f2c8f4b1",
      x"67df8c02b4a2ee17a8ce1f835840c72e7520d49b1196879429fac317138ebae4",
      x"9f57846494c37f699f7fcf14a1f028a015aa7627dbd566d02f89151acda38c02",
      x"be9f5ae493935dc644d7c4ec6910807dc462803b23f48b129ff1c057c2abb61f",
      x"8beb8a3217ccab60bedeeb71c99b81f5bf7c3c2074ccacf08fccebfc1c5f14c0",
      x"69886934f6e369fbbc43424ac614bd120c335ca13f70b00b57b7f5b1c778db42",
      x"dae075e9969450cfaba0b6e8a7f2c4428cb1fefa0e4e85b165c6070cfe8441fd",
      x"9d56d1628066234921541305e42a2a29c85a33d1a65be2ddc88f688acd4e2e61",
      x"2aa854a739e1c799a733f6323ecf163ba7241b4316a3e170c843974957f085e2",
      x"f282d4290385806a88a0d06db122e38abe46934089b13062ea4b817cbbbe443a",
      x"d00b0e0f0ad7c787f0d89edbeafceebde74fb863116db027484a57985db287d7",
      x"39b26c8402d1d81f92d16eed538c3ec2032393788da265389c52b44f0f86bff6",
      x"def3e2178a62a3bd6548fab949bd017b157aa5e5bfb18117162f8c47c9d16352",
      x"b0abc3ad707f8b0ceaa9941ed1390744a45253da71916c1a8e85dcb06f48198f",
      x"6e2aabc6b28e7e20cd854adc9e642c0a2f78f393de245e58a45d64c8c8ba1bbe",
      x"e70dcd5cf96947a133c47e09f3ce8834a8feb4cdc74c9c774a297a84bfc0f3df",
      x"16c4c201af1a199091ff9e85ddc01564c676f286c90cd5642c7debacbafe3408",
      x"c62406a45fab05d89014dccc66a9141dec58232deb84e4396a549922745fab18",
      x"87497a245226eb3a51bd38cb9d936f989bc74fce768ac67ad24f707999d92971",
      x"3fbc1fb40d30acf290f327de2ed2e5be01918f89e339abbbe31180178ac1ecdc",
      x"d68b297d8838fc59e0692f4b86673455d61f84db4141f109a1facbaa1cfdb367",
      x"047c03f8c0a5d1158a42efc29b314a9a6f4a5a42c9f20ab2c30ff8d45166a8bd",
      x"10540f04e26917255a126f599c2132c47a773c0bcdfe7e084a3f3e41711eba00",
      x"07bb71dec4d3add21e753fa2797909775e9cbfa2ec683d99587fc7d6e4dec9e7",
      x"a16de6325e6dc4f522e8f2de7409448aa4f180d1385696a9063081b74f44d4cf",
      x"cc5bd0ea378172fd8e0bd07c3030f30367a82ae7536b88b42d6bc9c00101168a",
      x"918051dc7e7d0c1bcbdecd0eab295b0461ac9b03374dc28553275718c6dcbe17",
      x"fdb67ab47107f2643a507c6fb1c4a71a8c4ce9c4e62ce518958b0b5470e9f70c",
      x"7b7088443701b3e80afc45f2e773f9d1c3ffc80399a639b55b5a102dd28d0387",
      x"4f340feb4062c898d078e4dfaa7e11039a0ef66efdcf014c7257e45bcde77c80",
      x"7d42f2649e1b0054541007501ddd6147a314ab5c126440df9d8e80e92167a434",
      x"b93aaaa7f90cde56600bdfd5bcdda421afb3afd751105ad9c1f587c7e3f70c33",
      x"4c9095dabe9a9a6cbd2dfe1b769a6553a92241104a66a05b1e24ad008b742cc5",
      x"bac2ab893bf41cad45faafeef941d8916e114ed5d4f34f365b30eb802097f29c",
      x"c88b8a271f625d3339b18963703b781c28123ffab1c4f57801f8706e4af6232e",
      x"331a2fe469ed6bda5a28912c7d549052776e7f219e22522a6437c7a4c4211ba1",
      x"037bad2ed49d87bc77b2399f63053f0bd6fb76c043726a33827e22d29952e3b7",
      x"6de7e1537e21e4adad083661e9b16f40087e4b09d8cb55080341a0ee158200fd",
      x"ee0ed5031c4cbc8d51d0b7f5201a070a1b3d754957223cd4d60e53164a3fee97",
      x"f41169e7eeb890dee23dd29d653e1f1527ea9ce77b594f752db07cf1b0c80ada",
      x"cfaa58412d49e720ca9c668341d0a239c592ccfe764976d7a746e0b4c372a781",
      x"b6e29d6172c264e76bde43ad0c332140ace15ba14464c9d81cca33aba2a895fc",
      x"bc2b08608295a8596088c02a3661d5236eb2fd71ff611a60f6095b2a6a9ea9aa",
      x"a5c132c39ef5385c2ee4ba34931314f7f1a45c634725323a8c37880254a15449",
      x"675478e8b73ca5f8f6148bf1817294e8f8764d2822b3f748802d476d07ddd990",
      x"c38b7b3cc67a97e66b2c48f1f97baf9f87d75e2b2873f0ef692325fb497386ee",
      x"19570461e0d8c1a6b2aebc9517788572e357b3c45fd0b860ed00580f85ebba50",
      x"5f5ab861d254a8af789c7f76efaffcb39ff8307a76863e05df76439772a19222",
      x"8b626481b5ab80bd84d7ca5fed1b9437b57dd951b754a9007fb73ff49925ec65",
      x"80ad66ece2c747690236404f45fea7f624a2f2e8f975813715b01892033352b6",
      x"c0e245ab7622ba616ecb39c1d67023012659c19a0bfde4cf5bfc9ba47608c473",
      x"9a9acd4aa7a334750c27e0a1801499ab9c68af6c5f6f4e1769fd5d1499fca941",
      x"d7027edb24c0a609361ad7beb188d68338bbc8c6a960fdb708d28e9ee8dfccae",
      x"80d6a7b405df42d09d30ab049cbf545b240132ae5ae28155f1cd683714c176ae",
      x"9b579ef9207a77ad5fb220c4669de18ac67fe7f54f229c9737bedff323324147",
      x"73f3e4b612bd2d76b08813751b79a113861afec9a773aa7e4c5152ace3d20e16",
      x"c78fec21a00bff8f05198552d400df778ae5d26b941521aff2bd510ec9ae0ff7",
      x"06fa7584f7b7110a5c9036956d7b0a2e42c004727c76c0b72b38fc8b2f64feec",
      x"72106053d8b956dd15ee72e1f387f13c686817cedf28cef357dd1a7594fdffc5",
      x"c11a8072e99d808ad2eeb1f412894b420279b84a95b4dc9554cfd9cc6856bb09",
      x"61316aed531e72d6e154f46ab3877369c3e0df14a01622a0997085a1f9229562",
      x"dcb33f16c65c2ac5f49b946c2f4dbf1c831554ef8e36e0bfe85e579217ea19bf",
      x"59701ea7be057bf27cc5e8aa1028a73348fc9cdc644375f80229979260134734",
      x"22a3c4ff520aac7da921d48e61fc6380b18392a26ddee38bfae29f587655124a",
      x"cdcf7cac57d62d8ab8084c900b7f34fb2d4f2d36126028fb7cdbb36fc6f38b64",
      x"448c13ea28cb8b099ebcfa3df26651652fd256971b4bf05a73aa7c866f1419f8",
      x"81e959cb47cd90d5959371c589b73aab4f48734f2de39929c17da923715422f7",
      x"0e527fc4f5fb1c50fff0d4cb7ae1086475ed1dbec6c564bc1aa2ef0933d820d5",
      x"7d6a954a49c5ac21491f12d317051c431fc6b330643bc829ed68e3f35ad24fc0",
      x"86756478e034d266ce3f190b00f95216bc0a7f2a1864fc1cc03d19457c6d44b8",
      x"1eda757c854e18e4d714cf8bd26c167ad29a29e800ada80371603421ec677735",
      x"888264266b0681297aaf741252472a0fed4ece67284774f2ac6775bb66f050eb",
      x"9ec104fa0c8daf9b7465e763a44ea4270e565d682910c2ad48c94d7df262b0d5",
      x"6cc2a675fa197c3bc51e0e77253146d57d42aa278e6a72e37a0d971027c96ad6",
      x"044347836c2bafb80e2377b77fe455afe1d674c04fb00258c982e5c4561bca17",
      x"8fc39f28a153e515b677ea1b3e40322242ff24960bc73924a011ddfaa285b190",
      x"12c9a54cbab7b0acf2a8dea518673360b9161d1767199d9b3c4c5306a0f0b214",
      x"41fc3bced33ea4c997a62d74cf0ed2d3cfad267035326ec8a5c7f466ee63b14e",
      x"4d957afd8f57001bf20694429162015d75557283b1d99bd7a9ece6a2b201ccf9",
      x"508571dc67568f7afba474d4df2c7a5f6303e54dfeacc3f1c1aee0aab0ec3424",
      x"2f08ebe535686fa3faf9f0c38770df0e3b994aa7e18743a35bc68aa2855c7221",
      x"5533ae2834d732ca485e2a85f94b4ba2c8d844f1a1c152f473f59ff7457ead0c",
      x"545c633ebe8205c8c5c5e0a6021af370b0a6ee9293008e1854f8c87080079e7b",
      x"e0528f24dc99eb30eb014d9064d0aad3d44a92340046c7c39c4612bd53277585",
      x"e4f20917e92be6ac6eba926cee4ef591ba59f87d22093828b59374cddc7ebea2",
      x"a8eafd7d00e0ec592b9730baa162387cbae606767cca980061237f84741dba8a",
      x"6205bb0ed90bcf2e20763cfec26e3af4eac7d5afe20a9a22ee26dca1a456a01d",
      x"3504fa056a043f1d770aeec184576d58798f0218ffc36b93232a07d27d4a7a2b",
      x"5ddbf9330a4b674926399ca44816ead0c6097f2d6c42ac0eb78f9e717bf0b98d",
      x"bf2551d32a2aeeb22a2fe4c2d1020a3ea41b60132d8207073425f87969b56656",
      x"08deca0afeafd801ebc4f76b00ccba805d162e9d1704dda689eda5cdcd34bf03",
      x"8ff89e68323fbdaf01ac61ee186c9bc0d9e4eed56e18cbae429649d1fc1945c0",
      x"3b11716210564153f5cf8ad115ad74d75e2e1c70c9318280cc6303458aacf674",
      x"3eee1848ca1b63c0779b5e3f86997781e4aa2dd7edbd1a6dedf506c97dd22da8",
      x"bac34221c9f00c4bc326888ce251310aa8f5e63e33fd6fa68b9055e60804d777",
      x"c046cba27118199f94964be29237b9b104c55f4fd5a63b8b44c6ff489e5528cc",
      x"1fa995b6d173dc1c104582ed53e697e125b426731d4ef1952fc346704abb7f06",
      x"00fdd33787b89ab1b4a629d135589f93c2e42e71d907860a0fa8d423ca009c8d",
      x"b1ba18366eefc0cf2d6bfdf890c0d0ba2f32a8cecc645dbc0e7bae0c43acb053",
      x"a0ac4e5b89e6567afc912a8f6f158d09b8b9d66119e69b1a063d7c348df41014",
      x"7a2f0493ece4249b9a12099aa568854d6a174bcc0fe8b0f8a76ad16a851d9cc0",
      x"b83ac3c7848c38da08910b77dd07168865171b3be6241803c9537f85010563cb",
      x"b1537bf7e7b2a5fdc1cbda3c04f048bfcd602d1af36cee42f5b8603bc61de56b",
      x"6c24a4ae866e06e8b0e55db130cdb5fbc6919b90ec7b271c8d41de4f839aefd8",
      x"76c25e93d88f548c4d9dcf0e5e3003d11ac770711f92b1bd5598e93931132375",
      x"c302fbca96875868c70ec70b7e3801827ae1e1e29f590fef3ae51b4d405240ef",
      x"7feeaf5c336d235ca64aae176efaa3887e26dc1adbb3fdcd7ff4ff7672b9dfdf"
    ),
    (
      x"27b6cb93b6f860a4a74e3101480f15f26fecb12879a7d00b970fd553ad5b1e90",
      x"b0686cd11cc1b95bf6b6c5f2c98ed60be7c5eebff96df1abcf0c746fcc56a375",
      x"578333ec70896449ec42be9e1f0126b179a35f2314090b0b2364d98b2fcc7ca9",
      x"21d763cf86d3803a1765501537f0ee1cf21441587738835b867e98f6d3d91059",
      x"622d404887b87ec4192a18899efa22c49970aa41aaa6a4b840032aaa4f4745e8",
      x"b335a000ff2f3e77957346a20f9381bd9468c76c632fa2235c3c84ce685ee302",
      x"cdf67d4376aadcd5ece17d2b8ff57b03556e31029649e4fb9a5593f2965c011d",
      x"7a2a02f35917f0803902f07b3180f377d6188204ea68ff51682ec1ede938d4df",
      x"8c36622a016934a8ecf980b717d910f14ad59e2126a4c636d7cdac9b542d5ba9",
      x"b53980c162e873cc1523a3d2f91871aa973f115864707b34cd4d82e9be81d70e",
      x"7fc8da14807ea689ed5bd980fadeb20a07e1d3dde868d14fd7a65170aca6e2e1",
      x"4581c5e6c2adfb0e63b80f612a93b9c64656dd5bd6c221a43d6c3fd3ec3216f1",
      x"c0fc32aee6d16e62d5e0455546d5a4d23989bcf4a01706e9415d96517e16bcd8",
      x"2e50f89c0f9139435b60a7f1cd8d7138f5e35dc40d5a406d56638225b151c9ee",
      x"386a534be1df43578b938db0e9bae9ffc0372c9d7ecde7a541638309ffe1afe3",
      x"d7c35f3c6686d0f82298e9607e8cc8a6bf4b447fdd0bb6041c17132fb4bdf22b",
      x"96a31bc881c8c6c315a7e1dfd79c577e5c426c5ef2cf96209d5931291f60ae72",
      x"1bb54540bc563ac3ddf1c1722f3e7d47ce9827d0ba00952b4995487d78b98ca9",
      x"b5b5f2d90eea42e79924c4b237d4986e547eafd76f14cb6de223b5d9033f406c",
      x"16083d00ea5a65f317a694e6ccfeb3f2f1b5b6a8727615ecf016b8118309c937",
      x"843de9ab7c7431cd9ee53d2795d593aa2de26b6902e0187fe66453510911fd6c",
      x"1be5865c95fffe5aab5cc427d24dfcca7387a8310ff9f3d9e83d21a26ce90331",
      x"ec8509fd3bd6bf8c771e3a3c8e328bbdfe02157cfa939f6aa869a4a7c658d000",
      x"a9051a688c0ce0cfd99b3f317031fd63d76aac9f1bcf1b8c2d15a1cf44c45fdb",
      x"958c94865258bfe4e26561743f82e6ca79f4a7ef67b08fc8ee0871c7d30a96d7",
      x"9029e62fefadf4351f948bb75989c78b1d7cdf476f5f27446e1acc0e0e09d96e",
      x"ae3950e9e6fe7ec0b8627476ecbf26d6153901b061ac88ea5593e2fc7796df61",
      x"30f74587de63851cb6eafe0be0ec1069256dc142927cecd5629ed07f5312eaad",
      x"f2ce58363b2ea08f154014856743b22601605339dcbb90e0cb1e86f913e3aeea",
      x"fb45d9e329e4195032f45a19e27451e28c915aa9012f68c92ef31f264675f9a6",
      x"48eb7c8c7046d039e70f7c8076590294e1a25e999b9093b3c183b07bc668ddae",
      x"7711ee097f3c845e1d1d05c978a9675ab07aa54b75dda3bf8ebef5bf87ce41fc",
      x"c30024cf7d1e8bbed4257de0b9533e854b8b29f3289ccd667916307e6e911c55",
      x"cd8dca30dd13d1c6c8d0250abef501455b975c6048f9fcc059a0ba88d3a1b426",
      x"1bc362c0b5b746795f4c2d4ac72042134d79f385c2b818d36963edb21eaf436d",
      x"88f3fa36fe771180a6334ce6d7d016a590595fbc2138f1e6c5542f1888e2269a",
      x"3d72cb0bb113a14f22e32c3ac2964c5188490177f75c5b5d4e18af5f3e37b91a",
      x"90f269da40f113dd75da5e30a956bf0f7693b65d884b479ee809afb641d53887",
      x"0fa392872498591f488220c7a35c795fb4e6aa3571685be39ddffce48dcd0fb3",
      x"c0f05b1f0d638bace248651efd4378196d3b0eaba75a78ff63019f5f126bd554",
      x"93910869ceff9ce355cf9bcdb84d0030b1dd3c8c5a9b9682d49fa486e56aff9f",
      x"3b645cfa62ac5ea7e04afbc1d605f83f2fd9c4f2e9095318bcab1953a7852491",
      x"a718a0076522c0d74c1514f3b2eec1b17d2dde0545329405886cfad1f960d407",
      x"b219340bb687f3e3452c6b3f26e6599714500fd02fa2e00a8548d6e5273bc335",
      x"b9dda5477bded037b90a524ce92f30f2fe78e7e6275e57fbf31a904720b1fde7",
      x"65111cb0c988d0a6727be1e17f85f5034a867766fcd8ebb3012b37974f16a634",
      x"967403b8bac1e9b8cab92a8c5773141235de56e7f12798493c95910f528bf7bc",
      x"1d2eb4243d3b93b16bf45db400a14caf45d912072201689e84988f6433a8318f",
      x"f4fcfefe9a360805a6eec60b7034b99222bb6e9b7298db03e7e522c1960559dd",
      x"d986b4765b0fcbd809b42bf4132df6b3a3872b90d6c0a20914db6182f1220ddc",
      x"268c7700557c1cbc9f56ec2c697cb27ba0468ef73d1fa7fefb2da99472284d39",
      x"c7799cb6d6ab86e41d8e5e171f2e381684290d426dda2fab7304708fc5174b05",
      x"c0a0d8ccaf6fd598292cfaf92b0ab0e2308f6df7d395817824e11e290fbd4211",
      x"957a58b134eeb458388b6770bacf4cf28a878a0e3583554da434be5d085ce23e",
      x"02e1908237c458a692ae37abf5e25c0be885a5b95f2813bdbbb8300d995c2b5d",
      x"eb521dd5ebe3bb2d69149ad2e44726d377566ad4a28ca43e795e2fc713c420be",
      x"6beb6b0fb2922cf68e139773ce31eb69f1d60269d1daa3ac8436f8cc823658bc",
      x"f55daf2395b4bde7b5b1f8f7947ed14150b60b3480d3da7da02c5875683ba674",
      x"61b07bf2b0cde7cd169aaf869b50950680083c2c75a354a92a29089d7194606a",
      x"d27f78ffd8b4ab9da2b70ecae4b4ccafdfe6621671eabc2265e5633837c8ad20",
      x"352de037d25a3c1214940024736ab878e69f22f9ebfd2015f5a93bef6095ff1f",
      x"91ebe4a02f64ea3f4a3588b6b7836e7f5d6670b51a166485685bd51c1bac89a2",
      x"5f3617927ef0219bd74b353d00f96c8fe0291499107ed1c7e67e612448190a65",
      x"cd6d900d4debbcc6ef4528ce4c87e1ffb7e9ec0cdb2d48217911811de9e72ac2",
      x"c70de731534e855939398e14103b0cb0c0aef773dc49185207842b835399d756",
      x"b3189f99a5a849532387d0f64294553c27ddf22a57685264e0f6c1f8e3e4ff8c",
      x"fa7e43ba194cab1c1144fee0b36a92f40589efaeb44090cf5ec5d37a7a9d231d",
      x"fe095bff84d170b7ba0df26d1d99d8c6f62ecfa4ebd802c9beacfafa28fcca27",
      x"41e39de380eb70262699771db2fc8f30ded22d9196a4c65cbe34afa76b3dd950",
      x"75f88a89b5890bb677fbf9cdf3ae71d72bd3b7c5f5549ae03decd79de16852e8",
      x"c7b40c1948301b94481772f255d94d0c1b6ae4b82217fb4f93bfed97cbc0679c",
      x"c68339073fa0654edc75491e94f9acbb632cc90dff2b344cd35e6f30e3aabf5f",
      x"8248bacfdb983ec932a709bd6d758bdd92283f3361aeb7b216d78ff285a907f9",
      x"ff0442e2badf5195f98867288d5f197e0649ade5a82fa67f70e6886e8e2b9f14",
      x"02ee477d4278f8a714913438cfc7ea104ee565856b74439e3d957b6a57805a32",
      x"60d25427c0514be6931e1418989c8dbcdfd12f6bbf4b5febc4740585ea998733",
      x"0bb8e44d9b571404620bc1276b4d5871fddbf57253856570dd0183b01aed5c70",
      x"8217df0ab5c76015e2c6f9fc591b7f4c5af7eee2738c50b53aac45c06c127893",
      x"4d4a431cc8151fbab0f63daf1dea54c71f0b8a425ab38e090b13d829a71f0470",
      x"3b86758608fadb4747cddf1b2070f188b0550bd9e69cf40e71223ffbec8f367a",
      x"10a5ecb0dd46441f5779980d7d8d0576527751a88502be7138e308f3582382e7",
      x"081c5f13a3736942ac97eeff6eaf3cdb09a5e3a78d373d408ab71c37b2f70472",
      x"dc834d07771aa0d2e75eed0e7245ac8c3f68f2a1ebd3a952859ce2d39f92c68f",
      x"d5b297cb6f594447dc00df9defe26eabbafdf78031acd10d87cd01cb03d8638f",
      x"49a8fe1ad2b63d8e374dfe8f3da4bf513d92eedc0f6f7b4acff89bf48f1ad2ce",
      x"122b84a5862dd54651facdea7b3b782a460f60421bcde5b8de3bd0461cf05059",
      x"1c9b732f5ac21e40fd5a92ebcadc267060e976ecbd31f350383ea6057d383c1d",
      x"ab056b5c0d9792880e4a5cce99127f47e1b59610bba53a9b2fe4aff12cf25e5b",
      x"f0ab003425f774948ed84b18755da22d7f09bb631fd5f90c9cd4ccfcd7f5c0bb",
      x"893fd56b838710b88afd27529f31c20784555db18c9c2b33c37ecb631155980c",
      x"76dc8cecfafebd63a6c811fc6614787a769b714d46fc5e383f627453bdd6f543",
      x"783251b33630ee9b5639042a703db9adc05086b2696e69930c660eefc01b50de",
      x"95c24d1b5cfda3e695fffece56f758eebce1cbb22cd492168aab3fddf36ef33e",
      x"1e58d056bd29eaac814e49cbd47be32486a53c6152ee2ee6deef7806f628901f",
      x"ec44fedb7b3bace3c5b6a1b270c283792f50437dc7a8f11c8455e6bd08a613e9",
      x"7e2271d0d0530c51fd980ea0a136e202073207e5d8b9621940ca13071d7e4e10",
      x"470079dcb935781e20802c16ae316c99e855aa39a178d84a7cc9a9b45837c8f6",
      x"1e64e30c1f01d50307fbb1289efa3b45ee28c9969a4d1b1511d94a74543b9614",
      x"2165023055c1d5e5071691e786741b4c056f20d839a4dd5df1464ad6ca43b4fd",
      x"1d20ae94d1e9f83e83599f2712711f2a7f78916ed0a658e13bd545f0468fd35d",
      x"d50b0ea6e8dbf2af2763f5225fa8a4e27cddd488f784a9d57895224591006191",
      x"8de9e4b2971c8aa057ce4ba6c8f448ad4db1fcb1b0cbf53a961cc344622b758b",
      x"8bcc54db0ae3441534c7b0865ae995af1cf00d6a00da3e26b6c528cd4b641a32",
      x"7354ad799548f76a039895a8f6a5b8ca6b5aeacd5565f9675f284aa7ca5d68c7",
      x"3bf6ecacae6aebaae33b0b94026f6561ba67b3cb4bd2a18dccb426b221e7d9b1",
      x"e6493daaa7661828106d4f14a47e1be1ea550e8879f1e41241d157e804b20cc8",
      x"48f46433481163adad572cffadfb306411f4f19f177fbc559eb34478d413999f",
      x"3473541b7da65f2d0721fd371fb6045c32c58bff56f835fd330fc5f0b9fd6746",
      x"8c14bd0a7f3f5377d72ae09b4ecf86886fbdf125706f478b078597f623cb281c",
      x"2d26cc0c7c0c03e1fa323bb17ac34e030b959863b9b48d3456bc703cad400ef1",
      x"6785add4b8b346361f5f3b032ba9de2b7c1a3b33f563fab2793c64340a8e5d65",
      x"5e6c252b89cd4b3c15b2050fdb1ba50b53e9e676b05aa18a60a904cef707af75",
      x"c55a754445ad4fd9d8c025872c312c3e557904ddfc2de86daff6a1ecbfe72277",
      x"76037e920aaa38ad4f78983630c8478ba6a6fd6ac17584a2682cf7a9ea7bc5b3",
      x"e6287e0eeda20323bf37baccc53d3f5d3884c4c6c72059a4aa0cb352913209b8",
      x"c8635d8c5a2258d7f03c25a2c02bb6f7211c08f9736de0a2772f43d471797986",
      x"1d6c360e573b574bbd0a2fd2d9ebf14e1071521d7cc8265ee6ae2ed1c007d353",
      x"9da1edd5679919974a89dda1f3a1a165f53e3d39c56c4e26f325fd14e89c2649",
      x"278893a1dbbbdd42e34546d4a72176469ae1d0caa1e963166473f970b4851b17",
      x"dbce50e9a252ff6accbe511a0658f2b1c55b0bc032feedada7a2d6ce62e46478",
      x"2cc623be158404e18ff47c83d459505e3687ed3330062b3ed977d9be791718ec",
      x"7f4062a5c8a5c67b5c89f760812724bed450855225bea656020c3e52f8db29d8",
      x"a47a3e3066c1a38c2490b235c422604422e492fbfb52022b7c1d2b1f6982f09d",
      x"b81d61a1164b2f56421176eed4d2704e8d6f42f59d41868406baa9f68f7b8032",
      x"72e732ebba9b4ed210531346d592cfbc2c5318beaf383078030cdf5a985c56fa",
      x"3844c89ac70e044143485d1b9fde954105752f095dd0b78162588af0c57b9ee9",
      x"be611b715c91dbddf2188d673487cd1a7c38a24f14d29f061ff26d23e61c3804",
      x"54ab7fdaec6f4cd8fae0d3abbc49129673d284b171f6e28b1f47a9ed6be0658d",
      x"951c4b93151b3aea594375dc5290a7c2631f71e482e9edb41c587d422fe1dc94",
      x"22be6a4b01346053285f500f0a0f0688e73568cf0ca6212d4361a936e57658d1",
      x"0c761377d4d38dbdb376060dec090404f85a15c7bf6707151c672601426c1c0d",
      x"5a1ad792cc8cdf59dc75bd2dc7a3064d5d9e162d95f4c75a8caf84481a3391f8",
      x"ab7738e151d32d3589dd5ea9540a1ed35b529c75682ab109a1a24deb56c8cdf5",
      x"4925addf6a2795fc2c134d0c460aa2228080bde8720b8c9fb69e3daf17154367",
      x"2f0c8d4959d0906d2dba7a5bb645e99c930d06d6aa0386b9b39238f964bfc0be",
      x"f036995bb160b4ead3e88c50bb5bce509d42109a21cf6ec814b1b94eccbb718c",
      x"ff6412999499c4aa3ccfc24caee2ed7fe5e9379183b101b6ac7cc2c2d7310b9f",
      x"2b333e22a3548a8d97953fcc0801438a33d3b44e177873f27ecb52a6828def1b",
      x"9762d2413e746e257c59b7158424b5b0ce64c411e080cf78dbd865880539a767",
      x"5369faba728b6416061b49175c778b76fdee496029d868aa84ad2ba022297276",
      x"528273652dc27ccc53a9d940c0274c3c8de303015240a1260387a93892c4ce34",
      x"e89fcefee5fe9b97fa001ad92489990c74ab0776e07a3966c78010633620d37d",
      x"198e1b7945cd253ef46ce3c0c9624f2094f7956a4424f7d3e260c52ec0fe4c14",
      x"927f3cb0c442dc23611bb6f7da23e88b7357b5926990fcb460fd3f3b628f97c8",
      x"0b0b6f7975802ebf7bf6404e459ba660001d799cb91d93563382769e7b4dbd6b",
      x"6bd0639fc858e024bfb808581e555db3b009ed9bee4b8ea6e1501c6b7bd4bbf5",
      x"dc2a82d7de0c63b6879da3094a53b4755b103d25f90808cf0da5eeb1acb70f39",
      x"84fb1d6dcf94dd81dcd5533e03c83fb04ceb35a76e53ce860c3901a5ee562c76",
      x"e5bd3bfcee6219f1610e0b8fc8bf85c76213dcd510b6fd2c64be70fcc292fc1b",
      x"4f2782b85eb86c47963b2cbc8e01da350b95b4370248f74afd5ed009b28677dd",
      x"e9a5101ad432c818fce33592fe9b870cfdc23f0c6433d3708c43712d7d7ec481",
      x"41ebe68ea0ae95ecee4534f61c13a0d8851ea95bd04a53077d9d63543de21c64",
      x"561123f3229b578d9ba7b638b9ebc8d4ac1c5fd7f5a4789b136654a899cc9ec8",
      x"9d179854e872188b2422e8f108e70b6f3fed21756c9b614f31f5f24922311dba",
      x"879b24f3c804ec00e7694a7d3d1725142a45ad2f5a7ead8b5fddaaeaa14d767b",
      x"50d82088f1036481663e9f9b33f52f5ed2481b549be29c3ae79692ac94f4f429",
      x"cfe77420bcb74ae5df4d4d0c8fca17467a4bc32caf5e346389bae8979bef11b9",
      x"23c50971a3bb81d50a49ace6855fd853d2744253ad82af666a1421299199f630",
      x"c9f73243e53f97795ce1531641ccc3e9784878ab112e0105ec45e5605b0bb325",
      x"052a7c6692dabd7edee716d853ce2fe79bcbe2e92f3aa6a0822cacc7e30709ba",
      x"a2a661cef3b9d5dc570695ff200d534de3b279284f9faef45ca92346af805380",
      x"6787684877a04149eaf43ab97805c464910a76731254dc6d09f33ee20010b8c2",
      x"26345b3c9369bee55b4948011eef5ef5902c12af6f9d6e0ca7efe7b76d5dbf1d",
      x"f9eb029b98625f27e4ab0ccef7317d51ad269ad748c189dbd3b690aa267c3826",
      x"7c15d536702ad87eff5307ffcbe35effa7ac5866bd48094d392e6ee25905a3d3",
      x"0a4bd38d11bc69f1ea7f5f58639b5402db707b9184fc9438a77215b2afc366cc",
      x"79598d16d563487e798a3ee7cba214dfd06c54bb8c5dfe8359a2f7de88f17aef",
      x"cbae8e542029ca59214581bb50f85caa5ba43e265d22cb2b075aa0c4201babcf",
      x"65960970448cbbfc4f3143abb37f70e954819eb75532437467d74d045b02e3f2",
      x"f003969b79f59f0dfdbbeda349acd7276b8939dc2ffada221d1d48ba1462a699",
      x"8ec3994366b4334856577ab651c41be6f10c782060be17f12cdc99199befc043",
      x"48ec30e4d38bd7685378053391408c190428e814c765fc6375f36ab36518d542",
      x"bd979355d5764e740899a730315309c37f4a091a23c5350d2b005c659a4a70be",
      x"f3ac6469f6c7be77f8ef168c22c8ede4a6e0cfdc52e9950a96ce64c1b81fb2fb",
      x"e1decaee4d044199e6e4784b9bfdff6381ba9285e0b2ec418f464461c8f912fb",
      x"98d1ec6d47dc2f4d9423315daa12fa65a911125f3099721e1f4d0b331ad78e0b",
      x"4e170fad829eeefcb446315bae87e90a8745010809c6a82f105430ffd06a699e",
      x"b069d00f95e8757393eed81d741546faf584db7c5cf77532fc698b523cba2029",
      x"5af38432a7fca7bf424ea92805aff3b39c1d1128a3d598eea42862a399ce61d0",
      x"36d90dab62619d26d9c56c11225734500317a790455142a75eb9bbe4963f67ce",
      x"bbfc495c6a1d4bc14250d4f8423d2a282cbf5233776b61ca65bc624f86726be0",
      x"c815ecff84c1f069655c6166de452c2a9a8ab0060787fe5ab062ad740756c446",
      x"05d9f14eb486d55ae63509d184bd641c6efa6e9845dac157d021dc4de2828b13",
      x"05a728a6c3def4dcaa9327469b6eb80918feaacd3f461f49b906c2b3935dbc1a",
      x"7a523f2c1b0a4b7e06dfe27b37769093576d43da72fe38938d97e451778fb3cd",
      x"50aefd08481fb951b7666b128f64501ddf1950cdffc788d54504e3243327b4f6",
      x"566070aef1a1142e5c0579054192a8ef8e9b7f8599a3031d4ffcf5424f5a93b6",
      x"6d215688a53241e35f0e8c39de5c1f659b6bb1d187e8076f11c0e19d634599ab",
      x"27b3a3d2fe87cabdd2c0104a5a685de6489b8f3137f940d34348a18ffc77751f",
      x"53497eb4cb51c9ac7458b0a2bbcd5a2b024a38b71a9af55da0fb289caa1f1953",
      x"d59dae65675a4d076695362bed87d9d0b5f542cd0a99b72adefcff58a753e7c2",
      x"49431a8468980343183deafd15b20ae008fb4e3782f9a0fa9d810aa48dbad0ee",
      x"91784ce8da112eb19d7da390112ec52e9cd662564dedf16128a018cccde39b97",
      x"def71c2ba0d96364a8c017adbb7e6b6216ed8f8d75a6ddf205715fcde048b4f5",
      x"63aaaf7b9d7ed2ac1017b0751a83fd76f82217770dfffbaaa9ea6e0bedf57572",
      x"02d0c3429b199b687c155fd8c861ed006e3425b8bebf6002411a25eb04a135e4",
      x"e53991ae6bb169c7dff604fe5d05fc88e4670eee5837af794028f4e36b724c72",
      x"92eaf36ef2bf9426fd67518469ea21c9fd655a12cd8b6935c07c57fc56fc87ea",
      x"6de9f36fc0220477166976983b7de5cd66bec1b6854936f2632e3762e2602d87",
      x"f2336426e2e27cf67c2b3d9ccbc7fe42344e016dd586c57db745823156f01ad4",
      x"eabf44d4fc6cc02342f95ee921b7c1dd8124007110c6941c050adf4367e0eb4b",
      x"ff18c6efc3f66be33c923778ddf022fe0afc0a7499250aace323b9912fe26051",
      x"3cc4c930eb96142f918d8c618b6f2e2a622e08be970786a782ccb8d17c1eae2d",
      x"d912894c56d9b2e2d30e8932bebfb8203cfbbeadd26cbe1f7a3082922ea36fb3",
      x"7c8744d38d5c95e477be08436a366ccec207cfcc7df1032d71a611569f33795d",
      x"b57bf796aa93a75a1b9a44709c04b991f6d80bbbc4a2bb906f131c3868e97e13",
      x"e4fa1c7686aaeb554357014553f08c6e665abf1d6883a232502ec147fd83df31",
      x"4602c2e026962db8e53bc0e36e5c2e53a23a0c6f33a237c9327280cb8afb42f3",
      x"f2bdf0d68d4be12d4bf8fc0991c443cc56f3694bf0f4e4c50eb262842e2a2dcc",
      x"fa85d8908e742e108f54989ffdb67b368f2a85919902aad1734296e852128738",
      x"d511918ca896817caca7d025043398bdf089a641f8f2475a40255e4de7ba273d",
      x"35166b89d303a4b8eaeca5822a0360fff8fd257a397e66032b4763e64ad9a6c1",
      x"26cc4a32ed591ab88674c33654aba398880d0aa7fafbd79d0ad24017cbad4ebb",
      x"d1e0cbb176e3bda39f7d2548a5fb834e263790117eb3fbf5f21013877e37a8d8",
      x"8e99e9dccb4135ce95bb5d5a42ef9557570a9356d41c4fd2ba356d702f80dea0",
      x"9d831f709d014360e4a0726877b644708c224164ac89d9a23bcd3a3506ff2536",
      x"b846ebb31e73a309ccc5230bc5e73d7b58b405f142872cd426bdeda7e1aa5a20",
      x"c6707407988392fc9631f8d91d324bae5a691fbde8e1999f67cec25e27a26464",
      x"2bff950cb85a2ff263f80d228e58e6467f0bb068b8eade0f01c8a2bb326f4758",
      x"3544e6db55f0a84c8cc99dcfccba3397695d01dfd23eb6a09d7369849a055a31",
      x"94ca612602167305d81ab90a112539675972b18abe389c0c0fe649eb5ecdfe81",
      x"78878aee75819cff41ccafec56044381777e1365dc202ff152c3d149b1286721",
      x"3349286e249fdad337945aa13fa9f6f9feea3c2517616eefdfc8ef8fd23b8521",
      x"c44181789fd6788737b3ff8ef256c6e9c4da168cfde8f58f05e32ca6c4d40488",
      x"faf2a5901b50d36fd4b8a0c859d584a3ee63f1d5623597ad334e02a5c97e4ce8",
      x"c2aad8225f5bf43ae0ee54cf93e4759b36a6d5dd20b3b799511cea1998badc28",
      x"7086af8c1579023c9297597bd15754dbba435e3b9e16dffc94f449b7156eae54",
      x"359270071042c9818cf7f5f69aa2b8df70696ef0d2e4efb4b5bfff5d79ce7e81",
      x"ed0685f77fb1f404052637923f8bf48d81954b390434d27f3fe1eb3d74dbe631",
      x"de47687ebac4112530d05854dc730d660e3dbcf592d21b4ed8492cf82fc307c8",
      x"aaa4161328714a64d539cae66d690481edc2eb1af17c647fbce140b70baa169f",
      x"a5f5c5d7e827e3017a4ea7fa8c92589a7f6b44c3e6453af2487bb7033a7a0cc1",
      x"5b1a1f782de2514a8209165e55125fcfec6a3dac71e9bd0d7bfecbaceac43cfb",
      x"b62998daeff1bce38faf9eeae0883c8fac3aa9675308df69e1027fda316eaae8",
      x"a755ce17da24032e72c60e5a69bf25c79edd19949e76c1fb1dfa1fe636fd564b",
      x"b3654bb7a984d11b0b71e3fdd71b4b2551b25bd57feeb65fbecae7eaa8628fd3",
      x"42f4f74eda1da8de6e98808e9ac78bf5cb54b12ef2518a62f8a95cbd11734e60",
      x"1de18f658de948a4d22ee9a29a76c8483ff3c723064daa5e5c50a3a82565173f",
      x"a7f3f50d33d5e9dd4333c25c1189f319af621a97490d6682279ec5b08bd21151",
      x"ae3ad23c6f43a8c3548ad441fc4715020e83a639be5c6628f6605749b762628b",
      x"2efbbfecd3a2953244b896d9b1a1e0387fec2392ccac543582c0b28c562a3581",
      x"d7a41751861f7e3e56c1c8e0a1a5852858fc3107f64ff06076be1202895a28f8",
      x"08edc75b513b7b0da62a4450f15d1cee82ef7ef9c8074cf565ea6b7e316a7114",
      x"a37b50a50ebacae9fcc392b7b180b40ee4a300e192a525fc049179f92ea80ab7",
      x"0bc4b6c08fbc74ae1e82cfe022100eafb905804f0c92094efc7d80229ec36708",
      x"4635faf6147348749b84f0b9565bf99313c5d7acb0df664defd0768b8c1da136",
      x"b2bc420c21357df8e3ded9a34c66a8a030e3142fd49c52cc69edb683b9562750",
      x"a875794ff70b04d401505586221d7bb15aa19bd77cb6b2b5de191c72b3625237",
      x"290680ca25dd64d74be9680f9b0266425c2c5ecad284ca94cbb290d5a902fc31",
      x"19de7cf141d96240ab542e8f203b45dd5ed42460a43a2aeb6e06fe6700c2d7eb",
      x"b5d156a28ecdaf830a4bfa956dd65708cc60f5453bd25bd332c31a1a3da3ebd2",
      x"0d4aad7286dcb8fdd743aa9516c8527b70d77cdc01ec0c09b4a57ebd2ad2a198",
      x"0f45c22eb63ed4f6c705a12666385955c03c65317a34af305764dc2261ee129d",
      x"68d86c9a09af9eb7d47b07f0351251a965b1f37c37d9d4c8c13de734de2b2253",
      x"e40e1fbca8e7511756a901b33f31c1bc52b188eb4f51ad0e30b6fe2385058611",
      x"5101e09bada9a0f41ae79ba39607345885c9d5bdbdf6b5f608c910b244f96000"
    ),
    (
      x"8129b74bef7411237afb9fdd0ee664f1801e425c9a11a9ccd33e5d0a3450e7f7",
      x"cd0854152294038a7b5e2617708ed027543ccbf6d54300988362caeb5352f0b4",
      x"3db2cb7c928ca501d3919d09f032b76c57c1f825b9ba4986c239fd60cbf42ac9",
      x"5b4fcfb9b349092d61179650d2e9e3eaf83b2c52aec75646e4cf09f4d8c1464e",
      x"92ab0e06f2849ab31779a860efafd67980dbee42ce6c5874e408bd744d3cb7f7",
      x"7612470200a410d10f5d0c1e7f18b90b5016efc311090fd720af5851f0884947",
      x"ce31d38578f3f00b12b697e4b716ededea11de09e487ed50bd487f0d076e2122",
      x"240ffa6892f9d6580297cd092728177a59d45295a403c0b4eb5a35120d604a5b",
      x"e55d4ec0279726d35137d0cbb42c5a03feb56fb4fec443b710a4a6941bd91811",
      x"d720aac6d500ae85d787251d0c84e749600df83fc8cc2398263249bd24526598",
      x"13d2f009dd0c3b516d0e652f58f0ec7eb04d5c624bda5cf6d13c415669e28d2e",
      x"77dae217a565a76ea280af9cd11605795819c6e38cde7eb9142f3ee013f78a69",
      x"f07a5a702afe480606bb88c2bad58d4db951eb170447a83be91f55c0eb5c898f",
      x"82f52373c58c6fe4e64ee2e33237c49a783c8ff8df4e55dce8bc989f8a9351d4",
      x"f16be40f82f6e3a96d6434816b1236576a50503e19149add07a0442c6f1bf823",
      x"0f8178e57bc7485924b259448529a0b42be2a6c0bc704a3bdbc6d4fcd99011f9",
      x"209913819241174bf107684d7ab1007e5150163a32e7deb060cb067ece2db270",
      x"22cbac145fe171e90b3cbb00485b51d975837d5cca5cd0c341a6cbc31f8c51f2",
      x"63eefdadce4f0c80ddd4aff1bd81d70b6c2d85f710a8eb141d3b712c9765ef27",
      x"a17d9af034ac9cef18954b798e587806a844396465319e5e34712f23d3c3e063",
      x"ff87d049b82fe5515f4f52f8d3f966b30b8d6db7493ec4d0b23c1b6cee20d16a",
      x"f3aa5e99b09cb752e51dd8a2ae23edea1e181a555df0ee3605d467fd1720281e",
      x"1c37a870766318fdc8ee120416437bd98b3c1126bfc28eab297fa5d933d6b0eb",
      x"85847c3ecce2fba24ec4279f864f0446072e5457f3d6d7490248f27f2816f154",
      x"4b04fbcb1b700d4a6b29f2aec4c5198533721b06aec9da99d86b25cee965ba00",
      x"6fbb1af516476b96ddfa2fb3bed30ff466cc49cc58047f5920711c5683e13407",
      x"a47a27ceb7a787eaadf8e9053a6df6c1f682a90b3914f17d9032caaa642ca55a",
      x"56d9b8195bcffec76f9b498dcd27a3413692344b811cccfa33b4c1eb4141e903",
      x"c6444ebc49917e85f5a44b310579ad65e8d23bf60d946183e0b0c722bc69da2a",
      x"b130ca0b8b1c789eaad4e69e7f54918735cc68bfb0219b527784989db6d44973",
      x"ad342a50981dc15624bb74733390d9aace091ba4f175ba00a3cb9e2952e55357",
      x"4556d8e6b5a012d69b7e0010fb47c1cedc53af971c44ecf2696447ebecbf534d",
      x"842f62100bf4b15221c25e578e14b249bf30c0579a51e0a9e7814604c539e37f",
      x"edd9fba566480b870586ae412a3862548378b22c84f1f447088f9de2383ec72b",
      x"99a6065258b9a6080bfa051f41797340b1c80024c1ba43e6946f7c1496855175",
      x"de321b32c4e634fcda982916c2319d21ea960f1baba36f8425fbadafc4b01c5a",
      x"43ae4e3d622576e26943a77e7b6d29009c0a7e1b0209427ddae9b2e3fdea1986",
      x"5a20897cc3af32f7d0b17ad9654cff72c7e90182eaa22f69afad93c4d7aa69ce",
      x"5a973c9083ad2ce1ad239b5976f8a21dffc64aed0162e55d9e101469e2300b34",
      x"89a51fd0ae44a701a8944bcce317a4b1264f5eb335fc313b67dd524c42d70505",
      x"835984e167b891392ca2d93de9f826699c0277e85953e0d62d2bd4594323da8c",
      x"c8ce52d56a879cb662134631b57d37090fb13a417cec36195f510d23526c54b9",
      x"6dc8da8f3abc909049bab9a5d8c78a7246a6545fd01edbb41372123d4818a24d",
      x"4cb4a92a79f562405cb6b6a12f66155021d02f9b22948440308f25668a2e3056",
      x"d5ed6429b0abd88e941028b5b3c6ef7c54cf72544a70b4703e929afb49596219",
      x"9a318befb18228575b5b421283d96a99c4212c64e8d3287a5c979dbed862e202",
      x"7fbc0eb27ccb47ae475fd6611d205c276dde1b564d8202051a9387f4bb81b399",
      x"1143c7d59ff761671bb065e09f11f55c4abcd4c77f8fdff53ad858af7bd0b332",
      x"0cad940e77b4bc8fcc3d0984f981c411f9a5f64126210b1054b669762bdccc01",
      x"128367726ef320f1e2942062265c607dd93c2f6ca242c2ba0722945da29c0593",
      x"2ece493924651a25cc7e91c364bea07ab5b73e4db34153ea8cdf0ae49661825d",
      x"f06749ca446b904bd1563f211be0fa8075018ef3b4170e85ee27ec7f94c13d8a",
      x"4a3fc99e37af855d11f393504cc67c2fb7c89cb5bdc55c6ae5d3a91f795d8e65",
      x"fb9d1738e457785147095d84250094e8788678e91d383a42b192b7b65101bafe",
      x"1c2933d55e2300bfe813787d61a1c30a7c778776bab589d12678a63bf4f438b2",
      x"0cdddf9097484762a371f5d894a2100426d212246cd00ac8aa15b47962c277a9",
      x"b41f0dece52390a5490ee16c7852d04c2ada2f0a778fd874f6ee3eaa57265ad8",
      x"02d5b975bd3428b3a15f67ff468f9e9c4e7a7374cc63fe6c99f13e1f346d0304",
      x"114c84d88bbd88c9903864bfc5b4a497b77e1861f8827d6dc82dc0b34ca72c00",
      x"5246977e3d29c34cc2e2b5739b72813e008c852e93631bc688cbeb2662b4e088",
      x"bc926ff297ff38b7d6a43e8b12a5f9708aeaf21272172815fd72831d77189159",
      x"e736398e9dbc19aa43e690e7db0794b3ebd4295a40958c005790e68e21a63443",
      x"9e1d7d81662171c1469ade2665ed09c9e52b290cd4777fd1d57367d77f65776e",
      x"59040f95a862ef074070873bab23733b2d01e35ba7798b0bfc9e64eed6d0b860",
      x"10ab610f48aa15bf361829f67d879bf7a578bc2a13dc40e9486e1a9aa92e7498",
      x"593628d063f101d6102198e8e547aaf3472021743592e95dda58bb46166ce618",
      x"7d9f992670f63465e0b9125876075986add614940dd92fbae43010029e775f89",
      x"829f47a93334b7089bfae5d58682bb698aceb851360667fe3a585ff7690e3a09",
      x"a0c57ec8ae010a0ead3e2243f5ef37df0598fc885349a625a03948b62e3e4678",
      x"ec1f9e6ad61751b00f3c11b1e9af7daf4f695e0ff2f7c193c353c74969b767da",
      x"330f427785686ea2135448909ecbadcb1dec62dc181bb4d17f4a06c4f9c3a968",
      x"6f17d585147adeb3dc0c56f0343c5d5e41305926ad3b519d5a9eacef0367c206",
      x"9ff34914084e9f415e2960d62f06b03c46f9e496710dd35fad2884eab144eee3",
      x"d1b158657a9da8b02f1938254de6f4b35aee5ef05146532750e0aca2fedc33b0",
      x"7f959605da7bee8141cbe53269cd3f38f6971ee74715812d9591fcc232ec1dab",
      x"b527a181a91ac4da5c615098e4b188c5a6b29631075a5b485a542a7b024de589",
      x"2078ce89f40515636d57cc72977aa2f38fdc55b131a9aa2b482c34836241fcea",
      x"227e4e8d809fa14319384e8daf1052ca22a1a3e4ad3cd0733d2e6ff538cbe5ad",
      x"a7b48af38bcec257fb7fdd90bf652664d30660fdd49992231d015dc8714262a4",
      x"1f368a5147d9400fce0ea863dc76eca0ec94db88fb1070f76847396a2c1930c2",
      x"d5dcf2267d95334de5e6ad326cb77ce5328cec7625fdbaf35d0a20043851da9a",
      x"55ec9e6f58a523d3582d07d721129908de3e44edfbddb0f4929c7aacb5c6d51b",
      x"5e090cce0f81dedba981375a9036d8a0f384012994eaa10f8a900b2398e29105",
      x"c099c517254d43cb8710476ed4758909afa5d9be1b498953816c75158d4a89a9",
      x"3ee1a3ede366bc96c8df0028860776d6e62ef51cbf1709053de1753e712e736c",
      x"b82aec9257313d7ccb55f226b624f72ab9b094bf37389073a1dc7474b4d23a34",
      x"1e9696f8821465cacd5d29e90c3fc38f4297c50677d6953d04bf3978a7108a44",
      x"4be925064d7d30336aafe029614d826581db8c6b67ae3c4b8f1c24ede08da881",
      x"d053e5ab52eafb600fb1cd6f5603ab01fba26eba726ef97b811235cc89ea2e7d",
      x"4d8a51b45fda54e2a4d202d1d58588aecbe000829631732fe6e81c1f4099dbbc",
      x"61b363c63fff9cc743ccb08bafc438ab7e41c4ed31bf52fd20f3face77ff4a3c",
      x"4bfb1cc46c41cfdfa9aa13f0fd755619ff9baf350202efe3b80b225910e560b9",
      x"4fede9660563abfcfd0d51900fab9041999705ffbced65df12419e6e21bb0bc9",
      x"ae2fe46d0734bc7c6c3e00073bb64c4a1714975bb12d1574bd646dded47501c6",
      x"a0df04fedacde5526311b16f5267eb17d7d024af3cb3685859ba2a6f149f18a9",
      x"083fff97c0f1db0600db2bd1420d4add750638684afc0b1324445c317051db14",
      x"44b6eff1add03dd42068173c1291afd39a35fc29d5628b31e2ee79b55a6dcdc0",
      x"4afa7137f32fe1d07ccefa77a9222e230b08e62d4adcbdb5dd8a2c1449f27b5b",
      x"3075649f8fbf1531ecc56c2d19f0b4de92503ee55af032cef557f41a3bdc0be2",
      x"98a67872938cb4f9713976afc0574077a35c8895bb7123a0f924ceb1c86c8e58",
      x"5b2debf5bdd9659c80c910b30f9ca660771e1fb3102d2e66ec704527aea9921d",
      x"b59ad77997c24df983ae6c597aa0d119fb907d804ff392fb921f2699252cb8a1",
      x"fd31be79c75576bfce441bfbec59aa136263b3dee3d0323f222ab8fb15a5f1ee",
      x"d9d32f9d59ae9fb4fb5384dcbe4c2465648500f81d7683d03a1be6e03d22f864",
      x"cabdb1d464c0a740ad0326a726629521076de08f07e9f632329f5bac773fc5a6",
      x"5aae7c25a21ddbb539460778662433c2986eeeddcce4a54a448d3451feb64187",
      x"fb478b4fdaef78821fb69d8492edb76dd5db86a55f08f9bd0b7eaf2ef61c373c",
      x"2928bb280a1f858cd5e99d2032e082cca4f19016498f7d9a8b4737c2361ff04b",
      x"e35abc24b07cb5ae0db0a1d2f373bf7461287e767a126096755a5f2cf1f3427b",
      x"99848ddf36113aaf229972532ab6d0f1e094a7379ea8543d85bd278d29857465",
      x"9f5e2e18c7fcdfbe87679a02be3ef970f0a440974efecdac76b08a2732b4a829",
      x"b7f1b8f8c5320599c9c4887e791be32d23792cfd9436f46ef2e05816f511d28f",
      x"1fee498a92e2edee43edc571607506b78e5a5167fe9ae8589a94b63b532d4a7a",
      x"9efa17f644710d6da8febf341c0bc3dd6c8b9dc3fd453ed42bb6f34ad56ee213",
      x"f897dade576fde2d93753f36729a79512bae1ab0d17fad795308a7c26dc5fe56",
      x"68fa3ab8da0a7160ef7ae2e56c990a865f741e6c3859eceb081f0f20a03882c4",
      x"2de581293d6cc5c8260ded1e84e9b89a0f71ea9adf259f633ef7dc36264cf88e",
      x"c3c5a6ef422120c3ae2a414ed346a7eeafbd53d9ebdbc8112d17260cb55df1ef",
      x"234bdb9fe05438f47670139bac93095ff045d31861b20484a82e717ce87e3f26",
      x"a7c9bfe7afe649de86decbf822ae4362c0bd1f26640ac449e8486a607ba43ae6",
      x"696bc7ebbef46b8d4df7038243b4bf01835d902ee1b5591d503823266ffe7e1b",
      x"556f49d24cb17a7210f060e61cbfd1afc56f03b8ded4f45f510c15cfc9d1edd8",
      x"4abe17155c5c145f5f041099b4464b492c5adbd7cbc24b98268420aab865ee03",
      x"67d2c517b862f3cb28cffafcaf965163d55af7e828c8ec963d09a639c49f4afa",
      x"de66887347657d1c0f314d8f34daa575bd376e97af2d74fb8d346e810988f80d",
      x"f38ccaf56858d0e22e826a8d9dc58dd29a5dc3d81afdcc5d0eb236bb4fec49ec",
      x"e983f71ab46cee00150f9c4328fa24ab27eee3bfa2fef7fe0d88acb749f7be7c",
      x"6c59c74b20bdd5064149b734b2ad2b6580d7a07a3b9fa7aba1b1a069e961263d",
      x"04778c7e7b44c8f7e0b39f4f987967fd382f59e23480eb1e9ac09209bca554f4",
      x"4331245041ba51df0e6523903109dfcf784d491670dffc5878438bd1911c183c",
      x"3da081631daaa99118121c51942850220a35d609c13f61ed278d827cdd83d112",
      x"ddcde2e38c85c8ab96f6f21ef19a696ac84b39406ebbefb4bb0b23b7f2a28cc6",
      x"5a76126163b912e15640dea3c496139ad33178bbfe188ae643695cb970cd3035",
      x"38391e74d7c647c324a55c10bc385a533bf1eeea45f7de51823496baccca774c",
      x"397eff9dfbd51d95a334b08358efdb93b7c63e2ae946fd862bde9d55e677b226",
      x"74da9ac7ef8c28e43f39defa87eba71dc0b3ba9272b8d1698f25e1ae13e92e3d",
      x"780b6a7c307f57b761f7e01d53d6cd3ea3daacca2c02757bca40ebfa6da4ea86",
      x"aaaec09bf20953ad0d7d2b12c0512fd2c732962eeaa81dc949c8757ab9140ae7",
      x"a16e7773312bc8827cc748c539cc964a134e9371a9258ee96d38552efa9f3da3",
      x"ccd988e8512912593965580cabced8ad544fd05ccc51139f86d777f28918d4e3",
      x"75d440ac2700511e75f9965ff7e2da93063201ea67e83eaad367c2b2218b824e",
      x"f226c600629d56addfa6a22af8e9c27dec17bfb6e7f705853754ed6e1db5501f",
      x"b405c2d720de76122af060c53c6504dd8040a92f687ce441d1c03e54833c2c54",
      x"0bb56fdb27b32280b74bffd24a74b6619f8c835a5fa56fd4d11ba5b7ebc9a652",
      x"6c1fb713d8a5ef25da9c7e2c9ebf8e8424f48f98d801695d1e7892e68953e33b",
      x"9dd8daad9c6ba6bd8b25561789ee99eb5df0ee71a8f9cec83451b299ca2b7949",
      x"bfe0057148dab223599a0da1cc5a61d39f86668f4ce0bdfe4467067fb2f45c56",
      x"724ca6856fa154fde84aafed71699d2419876ba5fa2f38ac9d3ee0013602b7b5",
      x"3cdd55d1ee945ce4381cbe9f96dffdbc475597681aa735dc74db1b3caca6f3f0",
      x"35eb70466d44f8349080a9647589146e1fa8cf6e628fa85f46c10cd50602f48f",
      x"879e8ab95651b9296cea2344f993c0bad31902e13cc44b9fb4d8c70bc61cf47a",
      x"bbe2caa251032aeee42daa13774cbe3577be1587052d70bf33dd0b8dde86affa",
      x"61bf865fb3cf14e313d0e425bcfc70f0cbad513577789c920ae4ab4d59869aaa",
      x"2b3f34a938450fad8d6694e954b607e0294618a29f4d7f7932d25a40850e2ed8",
      x"8e9f8ff0fd028ebfec834de062e0216b08587fd1f40868aa962253f5f6e5c297",
      x"5eeef0b94cd4c54347ba909255fcd622404bea580cbd610d8f065f33bf3d9af8",
      x"3f0cafe9578f9d3918abfb00b64f67ec8c124d6d6e7ae72a25b9765f4ae580e6",
      x"dae81d42e2c56fa521c6e8b02b90c8be190c05a370c6f2cb92f7d180b5c946d4",
      x"f381fed54a64e5cc15864cd903c316695eda6db486287f19d9f7808b040204a2",
      x"dc663efa472dc6b56672ff65f4664265ff94646e675eec5d545838e4bdd3692f",
      x"c727cddfe25acccaab3fb8204bb9d3431f17ac1dda48e7f56eee0e1cc0fdf8b9",
      x"520d7716c7c8fdb2ca0e0d87a2bed3e0479bbea6faaa3c5470a12796de67d5ea",
      x"06c871efebe63423b12926b5aff385d7979780bc507b4b1b3d93911fa79bdc43",
      x"2d0b49891bc7883789821b8caf257c84cdb170f0eb952dd3aba875348b06d563",
      x"8ff412cc79239d41fb8c8ae39a015157ef4757c6cb58f95a39a303004f4ea5c4",
      x"6ff42a06dd569c1e95bec99707d100b471caa917650896ff2d1dcdae411f27e0",
      x"ed67bc543683da005123e7d531e2457a0453721ee0c43e9c2a6cfe2e62471984",
      x"bb6963836919606d9f059bc0c362e2292854b7548b6875f276719999501dada3",
      x"6d794c4ae6f5dcff26070f8587bcecad6f6d5d2600dbb2411e1d80d5600c3d8a",
      x"1d7b6d8b72fd2b0a82b55c4be511ff96804ac44092eecc8b99214f23dbeb46fc",
      x"9ab2837c089553f48905a75184ec19319fab4a1b102271d2cbde15492b3a22a8",
      x"0fcecc1b99b8abe9aa71c5e98b8d48fee515bd069e8d8c6300e3acc8d6af4205",
      x"b019d35d8e5272e3a29c7bd1360e8beb5fd7d8f3fcc42e63008c2daccf7badcd",
      x"ec6292148d93a58b6df7fd12fc2dbb2535d4a6bf50e862a166e101e15f59d436",
      x"0d9434543c8eb7f6963f9d88d1ebcc8a7ea89e31a0e8e54eb5c92554b82bf90c",
      x"605723126980131a17d73b451f46151e411fe21972a6576f6e0924504a2ccafd",
      x"6fdc7e62dc973ca829c0ca65fa718c4918e6981a41f654804a909daec290fa15",
      x"94efa9ab8dd98fb42007c1925049cce84cc87ac1e4cf0faf880761500eca8a58",
      x"4c25d14fcdaf8de4e66f3ede375ef1c9063f5b69971b497cf0036357d64c9ab8",
      x"c9a8ca6d2acdc8c0979605fbf535b3a1c077cbb9ea555401cf4f64618d1a2be1",
      x"6fc1e39c9d08df639fa28f911d14332e39614c929f8309948a911ee426117814",
      x"20c43c995adfc1d74dcd4e692ec4be16ecd697be5c1e992b1a47f2d3ea8a2eb5",
      x"3a89c204286d4d5d82edb02bc69007f486374c8fa30bb4b1399c03a1290b0f27",
      x"9cf686df708d10cb928ca434f6239857b7a12db77e104e920f730ee627b88e87",
      x"6cd7b4306b04160272952bbae5c9b486a8de28c2336f76713eeed1c26c45dc56",
      x"02e585bd0f9d406dd9c3c4829a840010cec27c547d645b8ce88f08277f494999",
      x"5d60e541d90a6c3af2b22e6f90047b5d88c3a7faaaf8aa7dcc7c55359826fbfd",
      x"18b8db2b49100573d4f54cdad5b4da04df003e0e9f32924cabecd7c028b2ad47",
      x"bbf3884b61ff632d12b90f0598f401b4d5372f6cea55a489e427c3a436435308",
      x"6f2f395e2670c25fefebb8b509079fd371733472d7f284ddd03a1f89d52c8357",
      x"86822973475a9775212578adaf1330ed34e9b17fb21ce0eb602b342dd736021d",
      x"52ef5d27ef687a9672ed9b0548f878e2f0cf236ff39a16a3c6d7bd6598cb9942",
      x"de4400d29914e1e66945680971464f5a5b42de163ed6ebeb92313719eb19b43b",
      x"dd3ad38e8cf43d8b0b11f998e6c200167664378dccd98478af469da55df9fdff",
      x"196214e42ba07b7099950ff8828cad35ca8916155ff58a1c9fb47daffa57fc13",
      x"3a4a80f83d18067ebfd059f52426baf843d6ac5024a5f4620fec0fb76e6b259c",
      x"e07b3995517fb1f2b64c783aa7e3bc6b85ce68cb7cdd802d4d35b72ca41e591d",
      x"444c7bee242f505e3bcb04a59da73fd08902f64f503da6017bfee943dc09c806",
      x"b23716de8accb836b296d9c40e6f8e47b3851ca06db039d9488bbbd647b1447a",
      x"fe5f3fcd4f890b6452da4a2e67afd4185145f0d8f6e7116ff402b1efeb4ba68a",
      x"1d859492ee4863448ac35cae7450e6b0dc93697715441b19d24ce0d75c4b78a5",
      x"4f0ab295dadf06d7380593eb8376def7640d68c3d69361820f52f4012856bfeb",
      x"0994ca5751b668a3ec14b7b4ec169b733753bf911c2a43e2f0af3cb199b2edf6",
      x"381a6da5302bba23c72e161483333ba8c5dec457b07942b07bf98eb80ae8d90c",
      x"0a1a5149a0b2d39cdd751bdde290a319f061bf47d0a944bc2fb1b66ebb873162",
      x"b53ad03c244812f850c8f0bbfd2ebcb45d75c54d425aec3df19e8cb308d695bf",
      x"99efd0e62134962460003557b498c540a9c38ad801caa83e0d2dfc672f4916f0",
      x"308b7d6826536f5f6440eb0d95402c6d0a9e2fb18c5016107f7572b29b986340",
      x"948a77541e710ed7c09c3557ad11fba465c848b06e5943bad0829eaa1c23c033",
      x"628e70ab0680c5091c0c638b97d006085cb4a38f7ba3b965df94b9270932a6cd",
      x"121e05156c492372a18afab3f9bd5248cd9f08b3447009f339fc9da5c8cda343",
      x"23655d505fc4a05440e84d0e375c2792a3e9cf72b87e42896c68a5af786c12c2",
      x"0cac2164e21e2744b99f82fe59c01eed9fbe90a45c47273eac59b4125ef22f7b",
      x"1fc349fad7fa39f02a7cf408b11818f123b8def2002372d7f5fa4dcf8a961651",
      x"f34de1bdbe38012a1058f354c53579a6617e66e0e25b340cac31fe53b1febe94",
      x"c632e703b034bf40080ace2f7baa009f7de484e4851ba5d730f9646dfdcfcb40",
      x"e19fedd5e0d0fbb851ba3e5603c6d38d96a6eeea571eceaa943159be157be4ce",
      x"04026e033fbc27be787c34da77df721f6e23aa256e4081b681b7e8673a3362cb",
      x"ab524e1a162bf4f40e2735b9dc945b53667a5d7d9b14901fc49c0a2f4f798ac8",
      x"d1109bbff82553cafca11af31ab1f97c68a102b2e4d6097cd8d4a9ca3413f791",
      x"143a1335dd107edf22eef64aa81c1f3f50677a9fa6deaa5db3dd0689eceb6c2a",
      x"39d73c5691c1558032d178494316b94e571471087b542f31ed46925b89a4c70f",
      x"03826fa36f322285c679c05911bc400dec329b35491b9c6d98d2c615bdd897bc",
      x"ab5ddf1ca6cda6c12f01d9299e7f2bc6e384490d1a100e2402443361ef785034",
      x"d9ae3884a79c5ef4ef5d156a08bec072b5046c31d77f886fae3fb3443d4a2e8e",
      x"bcae963410b55534a4529fee265e82f5d9cc690ea15ec9c4e65ab2965640531f",
      x"7c2ff1af801c23e9c72ecd1dd104334e111692b0a364d717a67dbb4b1ef855e9",
      x"70f39397b5f95905a7bd2cda5eb44e3842266967f2760b117eb0018128847927",
      x"aa025a96f8e1b5804f9d95feace4aee355b6b74f05edcaee7679dfdf89237f1a",
      x"8a7a0dd8e1cbb9e0850efd9e009f9935a03587f02105b5252963a7c560fd243c",
      x"ad2cb1bb282aac4ec0a0bceabdf3b6058a5f0dba88c5e87cefcd766e4eecfe8e",
      x"6c24d371b9b2cc89adaf91b3cee4394d3c1b48745bc12c109a223ac1fc687da6",
      x"6058abf16a687e66f8d0155cc23c1b42cf83ad15a341f5dff01fb6991fc901f9",
      x"b77dc9788c4f82a50e105966661f096b382657773da93f9e7e700052f63c72f5",
      x"c49e271e5d7e25d9a97e65aa51b1a5d92ff879639c4e5f06ca4c3678692140e2",
      x"e2f960547fa817ae9d0c41c83351c9222fccaf3103e36e05e004ba5f0955899f",
      x"3a69cc3ba53916a4a02ed40d644a3c3c712bbe689eee56b4aab6ff9bbc724f92",
      x"e4021a9322e3bfc11f4a7f98aa5b63af2efb912615a72583b51c48cd0cb22d89",
      x"17279d7f1df79ffe7a2927030470efbfe290e63b9f9e9281a7e505f05ad50b02",
      x"f491b4c50dcf8dda65d80a929767a3a5a801a9b90fbd98ad4d29c68b85e8abcf",
      x"198c7b53d03546aa7f10fdfb36fce34e4ecc860c40001a45b536ebede300758a",
      x"078f264b8adb552134f1940359191836c6b28b1bd9b4345b190f02e6c6810f1e",
      x"c559ccf747f48dd1894fa85a3df5606570fff4afade65c5de2dc40c869e98b14",
      x"82b1417faeb812902dd8e3f32be007ed84ecb290fc72a75cc557358ca28cb483",
      x"e06d637266b92ef5110bca6ed4311b5a914a66cda26981073fe93bed442b5768",
      x"933af04071c9c81ce0f4c3ffdf835a69e2e584d45fb5b8790983846c84265aee",
      x"572204ec68fd3a14bc45d4f46ac2c5848783e05433e316fdf7c93fc3b9480890",
      x"8d1d3fee889c551c6842ee555bdf2186e69b037b90757b7c9a9e05bdce0a3ebb",
      x"725848fba95fd8092d3b23054e43ab001fdf2a27bcff8a115f7d91ac14e1ecd2",
      x"a0a158d81d0f38f78d5b32be56fc2dc99dd964682b03b85fd666626408588f32",
      x"db06a2e9b80035a623e41b304d7d60b59e3e65259507c2acdc4e44f595595b7a",
      x"c4ff2ecbcaf0306965d907a2bc15adef642481d4d704467cd445d46e180fd7f9",
      x"ae191d0b3f11c3f5a2f39bd882667c6568f02c60cea0a5029eeff8064da2eee6",
      x"22b7ac2d4c3c079064bf05bd4f849a17e2467ecdf9d8c15b473967fa1a7a508a",
      x"ff91afe02a6b5783a526b37b512e5ecec528ec19835a959a026e5d036d1b5cca",
      x"0befcf91089a1d1c613818961664f6f4d6086a612749becd1c680f27e1be01d1"
    ),
    (
      x"b33a0daadc974b7b9aeb6afa0e823bf882b8a422bb93587fb192d379dc1a7f5f",
      x"fea353565f2a47f2ffd96193bed541fb1aef901a695a1f57446007e3e2b4f454",
      x"4b1c9cb0f64623c05be844389232bf707eee5e58b911eb77de667d79f7d31808",
      x"6dce3107d2c980dd267a8059387e1d2b71a2646a5675823db1368769b4cd9d58",
      x"b4c8819392ab57e51561632999b34fb3147bb72d5606315b0bf9591f531f9e29",
      x"e6d592923443b78e40ccee098dfdcf2db5b107dd3b93cefd521fafdeb83ee225",
      x"af63d2a964fe98490420d67e24b37afaab016980b092508d456026967e3f9d3c",
      x"20ccd876c4c75ff88c05aaea9d539f1b1542fa5e03c2aa4e4c91e5dda05319f7",
      x"4235e1e634af3763e4017cd5dc662257f68b46bf2653972419a5ef31028b6354",
      x"fcaceb75ac731953cc0cc7f6843f72f400f3882ca13e6cff5bf756a48ff42412",
      x"892649ed26482b4a14db1449762276d0a653d40e78169d7a7e89317ad1d1e287",
      x"9e684a1b2da3dc12d544f257b5208e91335ad2f874433033276e6cddd79dd87c",
      x"3cf7e3ceeb1a90529e474051541f59e348bb8454bdafe8f69acf203b2b92d2ac",
      x"223b7333e04ce3eb7947e2e54c7f73da44773ec58b2dcc78b45dbe1c76af6d0c",
      x"7200a73f8587f090146f225868bdf02c8ba3e47bb33722d44f307b8e8f5489f9",
      x"462fc61671886c52e9de77f5e0f93d007843192f71edb389bad734f8d1183b6e",
      x"e8dfc6e46e5a7d27ab54cc030d103a6c2393b4567adcd513f66025d5f4a85193",
      x"dfc61cc657a0dcad2fe729b5dd8318911acc73a120daaed417bab05b342da13a",
      x"00aa192b7fc7c91494728a83e539f1a54fe2d32bc33f14efd362e0c43829044d",
      x"c9082bd97c1f3dbc3197c0dc6c7d92138c92a8280c957c0a276def028cfc64cd",
      x"1aa41e29a2079710fb7f99ca55db075f7aa9bd0c437e8db9cc5fffec6d43bace",
      x"19758b858b56168beb957b06cee45ea65a98167a3ecd996f23901ebef568b73e",
      x"97b3a9a8bb1b830572daa71e19f88b0e9b8c28adbbf328fd8052a4ac7ce9cb7c",
      x"f561804a8352ff1da94b013b2500f6957194141dfa3ed321ec5b8451bf9cbbea",
      x"d9d1cc3bd603b1e28043eccee5b2f8d8634a76b5bee621ed2b0ed1e88167b47a",
      x"abcbc8897c668d67397f56d208a974c26314d6821ee60e8b551a5cbc85f18206",
      x"26e626d6685edef5ba87e9411512bc7f36ab4f18483d86ea3c8fb9e2c06d6fee",
      x"2287355a74ccde30977ced309a2b80a18e71444a06f93fdbd3114f0be946fd45",
      x"9960d5bde59fbab3161aba82d887c9310c373763f386ba070febbf35f98c71d6",
      x"ecf8226581e83cc86fa722fae630a0263ba0e4cb9d50bc78d266165456554dfb",
      x"0d3355fe5c44df59df20fe2da8462809cff27cf7031ede76d9552169467ea502",
      x"70ba85e5d78a4fa740b8d8dbe3783ff0a39baed620db804ddd3806bc27a65ac6",
      x"83ebd433caefcab0fe5a256f98090d9bd6f589cd0014821ba3f9a6920641e479",
      x"5f4211bc30ec36fd8c1355b15c34cd91dcd26a33dca3bba523852c667e9d3261",
      x"33e807e6429ac01119431e02dee29a8fb7fd67f2b39d47dd995a1d3db0f9d17f",
      x"d3575b530a294d88c541131526dd3e87076b2ffd3a0738033485df730c98a0df",
      x"4aebc38aba2936c2e184f403ddfca6eb5c61dde0fb58d4214e9879be544461d3",
      x"ca9a07be8e5053bf5dd2486bafa4402e94aab241a71ed47d38088d530dac1765",
      x"f2db86496938034edb7f8390b204ccb34d6fe0c9bef50c3a316ab09ae4ee7fc8",
      x"1f169fd8540261441443678dc9bf9afbece158cce41d6d27859db9b3a2caee8c",
      x"551221cd1b3c60b296999249e2fe0ea02700870d98b81e3f8a9bdf7a1c3a3084",
      x"e0dac837b3e904c7788fab2de05e5570586cee3b87b8a378684d8b9feb62c732",
      x"02705a59bcc783782fb71060a1dd7475005ad0de36eda2e43a468cb017a39043",
      x"903c51d11b22be0efa8107f43cbd02384164841a1b72744152e89613b4b0137f",
      x"730d4d096c5bf546803b6af8bd2070e80deb6f69e059b684e42168e1436fa716",
      x"81726ee0f14d9d84abd30aeee5f46a514ba19b5039c0af98e2471e858a77df9c",
      x"fdc76d60e3dd3ee14dd3c9747415f2098cfacccb7c6431fa3159fada08289b6a",
      x"8279608c4b578ba45c0808bdaab4653dbd2e9a4e9d3e69a2b8178e95dd082070",
      x"1e53ecf45e0050a4ac6813f3baac10a46b8c5ef4e2995967e29dc8532700aca1",
      x"e507ad1e63a69cd28fb0d0f7b89e263a677ed3282ec81309fce80a8fe3218267",
      x"3c6133a2ceb8f04ed422856502deefe3b57ba73a26c8763907d39a1a3080351b",
      x"e32ca83696738a9a10078942af554f43cfd7d19359fd8670a329443ba2e20554",
      x"f5f98573f88871e0ccb147ebd2cbdbcf590455c1dfa79a9638b5cea2cd0edf09",
      x"33652c6cc4f0ab837d5efa3e3e712680ba4d26f1d9206673c510825d2fd6c5b6",
      x"8ef85c9fd3fd18a4c3e44987560653a9aa03d465ae6b99a401a9c7378a43205d",
      x"01f29375abcc0b72e9d790022f6970abea948ef34bda45a27166299c070127fc",
      x"82f92663835876753ce7e74b561d63a89436c44cd61646d1b64d433f9343a8ba",
      x"37ccf699b938448e246127e486e5ad6fa944c0e6681d3b2c9a853cc3278650aa",
      x"45fecbf3aafb01b99192ff0c3db954ced4568cc63e244db9105167713ec37f54",
      x"fede151fb304f9b0222fbfff1acc79322c42d596a1fa002d9dbbba6fb97ffdbd",
      x"d696a0da7ef66ff403ecfc7e6eeeb7ba91b2a9752e91f98a3ef1e1f26e4cc1eb",
      x"cfc69a49343ddf7363af4ed9bf11d694a09175eb49a594197173805f11ee70b7",
      x"16be5d940bba2ef23c58d0b177855070d42caef9adc90545ef9707c9ce641a94",
      x"ec8a18411afedce84b66efb25db1fbb293333fb4424d7b70ea83c484215ebe34",
      x"38ef4b7dba4cdd5ab82cc9ad4fee3366176b219f6f6ba4a521a030d43125cdd5",
      x"b137ee1f82df8092f3c44eb3845c93f2bd26328d5e30ad125cdaf57b6eee6263",
      x"960c3e21202eda88e362747dac595024ea1424850551c067ac35725f33f2c1c7",
      x"38f496fb580d870e43128851896017df5fd38e98eb99034523db04fcac63910a",
      x"d8d626a5363167b52b4ae2144aeef9810cc70fb322fb48d7358c20af671c3f3c",
      x"abb91ba4788a7bb984f501d2bb13205e1e9aacfabaaed4fc19127be8cd92d7e4",
      x"7c392f7e7258e8d90a9e0938ec3d906bdc52ec691cee27984e4eb3445739cab4",
      x"da401a54463846943f4ae395578ee763b52ada9421632220c07924c569080af5",
      x"f0fc4b62dd6ada71ab77d8061bd818730e66e633d0928e84474b3855f6897d74",
      x"c52fe8391a84d2e7eb55a3d31b8dabfec2a7b8aeb37d85f221b4ff41a377b627",
      x"e1fae549f546ef8a6e6856421db0e425ad72531ed49726c08d91f9fd32831027",
      x"4ec03b0e42c5331801168a3257b11093ec393ea4463edda708cdef770346c3df",
      x"325ebe3d44049d2630e4792c8f952e02c20832bca0fe98755f4de74d762c066d",
      x"064c5a5e893b8132ef6b23a4c980f8b1f034d390bcff1a4c56cd3c0556170966",
      x"0a22f174a1281cbf9f37a470dc052976b45ed6db02ac326bfc13f4d8bfc67906",
      x"51da6e9b84d959ad7f3406cd2f998017d9d82c105bdfbaaf680210a0eb49afc5",
      x"3dac0e8946506afb8f3a0864697314d99168cd6a281e9e8e734738c48da6e949",
      x"3480c5eb1ef1f767d242d23b9365566c851156c2a34bd12cc2d26e83bcf05003",
      x"2ea01d909a1d9bf3e12ba667a3f10f382f626f1e35cb03e822f3c6d9056baa5a",
      x"cc275b5e96390217f8e3d8135a1d814acb6842cd39b0f83e6eee3eb6153cb34c",
      x"f62ddf98b16710458a9e1587ab8d105377c087ee9d1445610753b5f5f4586745",
      x"b0495c157ade1adfc5b8875cb920c493833715c77c6f1b1aa41b1834d32c7e12",
      x"2ed43089cf167ebb8caba0dd025ed5c648b86d0e8e2d73e452eb436e8e3aa77f",
      x"f0c429d0b9bddd758aa2f5467720b2b533216891d81b711ce11cc61ac483c6a0",
      x"227e1f9580e863491b0262fa3bc796f49e2a386ebcb44f6343a7efc339c2713d",
      x"a6925e902f75f74f195cee8c0c31eb8eced74ea243e4062c16980fd7fd284d7a",
      x"bcae7c2f4d88754baba9a381acc5c148628754a38e7e0673bbdebe2e8283563e",
      x"82ded2411eff83cef8cc66f7855f59132ad6f1f5491bce93702603f2fd4c99b4",
      x"6012bae01f5054a732aefb2487aab55f34e847cc8b36165871b73442d1b52e7c",
      x"95fe9ae040a1d483c43ed9cf2cc08d86db010129b3d289ff1d79cc49a4114ec9",
      x"20b1faf96a811057c003cf6c6b3133a1c5c881aad457144d424421ce0f1e7d8e",
      x"e3fea388e968cca2834d56c10e41040b9014552ec66d1f671b51d4d2f0a16c2d",
      x"633f0d5819e720f9824e0bc8ebb4129aa625203f11935ef7283f245962f201b7",
      x"f458382862b821e0e6b4f88a4e1e1d3ee1ea673e432794d2182278687940d035",
      x"4c7840d83d0cbd79a7aff1caa82c17296a89015903fbde1cc5f7a6db2f52c550",
      x"f1a259cef101d67ab29bf7d4f2a7d159d405d82589b47b27ec410a91eef0e240",
      x"c2c807fd08c781d213d50749abe4cfd2ca9667a7815fed0ead1b9d72deb3c16d",
      x"7524fd81dfd03c2d97622c03f622524d3843e87d8da677b709f56b81b6cd1b88",
      x"5c2f55306898ab6fac1e8ecac880d91e334e633cf0c3019aefe9fdddf89fff39",
      x"78d436d1de3da3b2d736620a740567d04da21288c478f4f5358e4bea98309101",
      x"159b36ac7ce9b71e44a7a9dddca841ab8b796fb0f9b92aac36c0225c9f714219",
      x"16dd0b28324ec300e860eaf432ad7107fd04626fa257ce04f0c1d48875ca7324",
      x"810ef6cb58d1316dba40ae8bb98040a7df9d4de22520f3a00db57c69200f30b2",
      x"f17dafe597a251f7c229aa85cdd077ab4ac9a83830512688c85e7ca0c322e235",
      x"0c0eddb3203bc66fa1ce674ef17253d39ac0031553e6a9bfa208e833c06e679f",
      x"14b8355410acc87a0f5374a40e7e66d310484799b01d5509fe619e2a1d12a3c5",
      x"523ef325bd340a0982fb4b6584406d3c0889d1d94100fd679dfb51096fa1f11c",
      x"c3a22252edd6d9a01a92b595f67cf887217f39f3fc04fa0d2db0a8fa4e416fee",
      x"7b1385084c58d1b9402df13a72081b1972478ec8dbc82c9f6c82410130a2b21c",
      x"425602e612e9e43ed42659fa0f2b00b546aa70040d4eacd0c50746e3f6ce9d69",
      x"ebed9e98bc1063aba6dbc860a1ebe34c7a9a6cdbabb44bf1e8f62da0df20b0e4",
      x"20ff01627340ac3a4da2fd44847169ee98d67d3f5c8524a6d53b2b4932cb3f1e",
      x"ce548d50a3448489be5ac600a1d6ca2fd36ecfbff6819283aee7c85e8edb90d5",
      x"ac9741bfc0321ad9a84016a77243bc893d1bb2a01b1f4acff5278531662e6960",
      x"896de7d51d4ca7bcf874e53b6b79d206c906658d2295741629b237988799fc24",
      x"359e869c3606c946591469214fea61a62a3f90be9fbaedcfad6563118c444ca5",
      x"964109cf428fd8ba3e4252cb81a4d67ec11e3cf786fae499d95296389f9aa183",
      x"b0fe92a12ab6d16f7b25832136e2d09f49f74e3c513752a120b8ece224ab0185",
      x"6cb567c404d52dede8c6f9fd7d81403c3c6b58a97c8d68a9208180353150f3df",
      x"c4c6a23c442bb89bb8474b91eb323837a6cc649583d1b31e7b20bd5539d84b54",
      x"99653dec3883625b490f5dbe5a90572bf49fbec40dca0c492caf604c64040048",
      x"3bd620d3ff1f4dad070a3784bf86fbdf2b74ba8c194d5d34ef992033e0823239",
      x"29a8f0de7f88666a56bc769770a5b6911ed147aebf8efcf2499b35a836d9b462",
      x"8c5f6d52308c28fc0663ee3468e87571b4447125389702801e9716901ee26265",
      x"11a98be67344871aac1fdf3fd4684632fbf774ee32c3695c7e4358cccd2451b1",
      x"d03ed05dc15b89cb254c50e7895b6a6d296ed330e0343b4f2247b7feee91a245",
      x"0a0b62c76c6473c93230a157f57d05f4e0d3ff67e7bc36e64c2917cbe7bb2dc2",
      x"b2477359ca9b5dce6d4aa55c6480b8264d7d7765208b12966e58c2787a50fed0",
      x"2642f494c96c9fbb9ea3c4aa97f310211baffb3c6a91f40dd855094816487930",
      x"c6913e0bb57e6b94013f35357ef118148b490dec123aaaec40944e2e3ebf33d3",
      x"8e3ed4446e861c610e50dd4cdf598fa0103bf99f6ac8d8de028c731872e6dd3a",
      x"3cd149e247c36fef98ab54efc0abac165cd8fdae66302802b19fc4275dbae448",
      x"658e5b1b0dcf40cb2b0dae94ae59eea4c78e0020320bf5accdb809b554a155b0",
      x"475a3f3f16b80b38e0882fef036bb7010ac5269d0209bc3b1052e0430dd0a4b7",
      x"29e963ae53bd9ed64a5d70dc18104dae106fa99613ce2cda21cb1d9af03e58fc",
      x"8a36c644751aea5aeca961c7f981fc9c89f50935d3929b1428a0b0b3507c22df",
      x"208067369e6fb2fe92fd3655ca804e6c33af4cb9a43ea41e9c6b595464e7726b",
      x"53ef128123524ee9938d202850e10214cb138072f417666af777e4058a15ff93",
      x"8dd52fe79c4c410ffb2a0676cd4c3ab6f8920f668c3ae7de62bcd1192b6e6622",
      x"93cca81a64ac3389097d0e94b6c9c47f2a8e5568d515bbb7fcb9d5ae8fdadd96",
      x"bc9605d1a8a5130f075376d3f5e7709f46d58c346e11376df7606374c5fd87eb",
      x"b007e3f9d317c7e2d6aa6ab547c5648449f4568bbccf2382e1af17a8a1fa27a0",
      x"9bc684f3682200116a2c4588eafd600f9a938bc97a6e79fd01c8e647b1b08c22",
      x"e983e2febf4e29d6c0f8af75914945b05df1171203ddbde0462939d189e01a6c",
      x"3c44a71533811fb018c94984a54c2de2bf39ea86e0d04c3fdf90cdb007485c91",
      x"d1d81a0ae450b511dfa677af6bcbaacb7ea7f4acaecefceb4ebea7885ece1fe6",
      x"017d04ae1110c03a408b7c83f8ac6041aef1bb7bb21679696f7b6e5dd13e62e1",
      x"e6a4ae61b15a68f4c7f76824fc6c6f5434d248082a53c4b86bd72e78fa5ab8b5",
      x"6f402499284291a9026decf3e3b9c10fc87b797131fb49ed52187d3f8347c3df",
      x"d2b5879f6951833030abb9fd24a63d31c7279d4776a0dcf9953ca36d0879e877",
      x"05fbafd7e0a6ac0519a547f6a7b075378281833f08a4bb7c2789c6ec78bf104b",
      x"c1463d32c058ed62b986fc7965bbaea8bfd6a6b01d7f6f4a518bf4b181c25db7",
      x"f453c25a62f6fa007381ee8b839ad6be84b279962b11a02d68b0654f02df6b9a",
      x"e923ee2e455c40c21f30bcf8e61f9d8205118987c8155e93dfdc26698e1c47c4",
      x"2ccfd711f04164c8c58a98005275672c9aa63543c2dfbb0e01da5751b6c8762d",
      x"0ce5caf1d29fedb40b2940986e41d4e131bcfffaba1c0dc4ec596c1f707abc45",
      x"f839c3ac40b7d68ea25174080a4c838a17a1738142bd8c122b206e813e39ca52",
      x"966eedc1ec7a9b4cedb0ab63de7136182dec35a4696959be161448e6970c48a6",
      x"190e5b615e483df550dd3e91d1baa32b3edd7c760555227722f63bb5bf7299a1",
      x"dc7e7ba6bfa9601d8f163ac5cbe4a4464930c03a4067d94809b0afba61118843",
      x"bdfbf18457e5ad5361dd32c440db8efdd629086b0fdbf83ff7f4682869b8fa82",
      x"b32a756935377cb80fe4e179c9344e1223886018def5e04c279b7b8387de2872",
      x"2dec5facfeae60165545c5f6061d075cce06067715d379107cf663b6a3ed6381",
      x"19407b94882179b40b5793a9d8e68f47e2787d0bffd3ce071db716f80d9a1d71",
      x"d7897bd160e0802f7aa298934ef771b9ecaf7f03146787e0f4f96723c91d0f29",
      x"fe133c8daad263946e3c04455761ee0ed3b3fc7022da29654e0baca5c1f47946",
      x"e1948acdeb6c4a681bd81fb2c82f44cd57f1ce15fd5e421b9c7bbe1259907029",
      x"3ed76dfb65927a1312059d6239bb4da69242ef20102526a461e512f39347ff02",
      x"cbd4457a3b55388a7ff63e52507ad903f0abc5860e246c0fe8e54355996bcf35",
      x"e6beb42492b1d9155d80630701cd128a7e08cdcd0ba215e7d707c8d091a1723b",
      x"20544c811d38c78f29d3957293b8a3526d68adf434c16a8ac36db014bf8ef40d",
      x"bf42684b7d5fb71e211f8bdba28311fe7f6f9edec331812095bdb4b2e4c9723f",
      x"c03ea7aefbb7ea7943362acbe7d4db099f0a8a3ae4f29878d66011b3c086f34f",
      x"3cee78e862cbf764573a87b686923d6276d9e2b12af1f3334be3d7f91f42350b",
      x"59a53f90a9b1d68a2b24b36aba51d5b679e7f8b7e717a0a033f066a0f17d2088",
      x"87f3c73f1c183041dfe9e522bb97ecc97e6df1cf4623d173b6129d37e4f50df2",
      x"01c79d2f5dab96094ee626f42eb7bdfda260f06021d7a6975996596bfdabe41f",
      x"445b083ddf02c6c838ae1e038ec1b757ba9c950adb863f99c03ebfdc926e1121",
      x"bb469efeec68f5534a3acabeb19e3ba4be7e39a6f24956bba8d6350cdcafe70f",
      x"ac2a6677dd10b98c39f1408234d1883b6de177e06f75bb29b39908d0e1c39551",
      x"6968fe43fad543a538099631ba17356d9494266c94962dba033ec9c88300306c",
      x"8a2cb128e2de5c3eeb1a33bd877b25454a694e5f9485e2c52f7fe2bae74efe58",
      x"397f4a91ff918259ec2521014300307d1e42310eb3a65042fb7127bb2441655b",
      x"1ab726f38639ff599ded27f83f63e74ce22f3c8bff4f95275dd3ad638b29782c",
      x"10aef43e5d034a7bcc5a8ba700d13a49c0463f365d87188c856ef4ffd6bd7c85",
      x"2944cc7b2165bdf9460f6a354f10267e43879ebe7e1aca8de22fca55e6172f36",
      x"c0634652029f9c649343e477ba81b27cf5f2c9dbb57691630292a21119a78dc3",
      x"4d502410ec11bd09112dcecaca866562d3310c518f7f63fe4a642c78411af611",
      x"9445f5bfba8bce86b7f6ce7d3aee88f19af061a76a95daa711227af0e7a29d68",
      x"77fc01261b85543ad7c62a2ebb864936ae43dbd650f8faa750dbb4fdcc36c11d",
      x"fd8a1823a4113811fc11246b4229e3482ff3bc20071e13a42405548b3e922564",
      x"776dd30a8dc6e92744f01918bc29f3169629b0d0c51479ac2294aa27815fbb06",
      x"8e54f9d5f623cb8a7797cb0618c653080dca65f23bdd07a37e44e09037558e48",
      x"a63af536df64aab079f7ce0220e9cac512ba435c5e7de6c763cd18a8d4a21db0",
      x"24c6ad688179a96e768aecc19b21002269f7db138f51dae830c06d4a70784ab6",
      x"c5b104b1a9410a861e9b98c0462fed5a0f0347f8ab76707b71206dc37d78e496",
      x"d040d63f64e18567dc313dc725bbb3ee528c9f7ba57adaf2ec4b2331d01e220b",
      x"44a58069cd7408ebe3734a901facde44bfb1035fad16384f133ada4c17baae48",
      x"6a57d2e7eb046fc15aed5fe8480aa0b14e495b51330f2d6c9ba4246be3c038e1",
      x"56514576b9d47188a5224fba0275b91d8dcc2f58f442758b136d3ebe7f197f30",
      x"cbd9710b9c5cf9dcca7b459f1435ce58cd73479f8307efddea24cee6fad600ee",
      x"7d6a1940f3bca29860fa75f8e0a1b5c6958d67916715db688f72e60dbb8ba76b",
      x"9ed7c71cb846b4310fa84a38e66e5ddb5e3fce83a4a4787771280637edb08939",
      x"3f3971401bc7ac0e2e91df12ebba304db25b5a6e63b35c012cf45fd51a4a8e8e",
      x"73e762bbc90e7e6714858b7f55dfb85e4e31cc212dc05a8a2460e5e3e5055d4c",
      x"a653e62b59d9d77d4236b2686addc69538e0c014195c823e3c62ced877f7ff61",
      x"ec25a3784dadc12042d3baad1043b03af96c4a6b133271adc14031c9b07504a0",
      x"188ef86236dbf3bf36816e5f5f76d980d991de2132ccb39b73bdf6c2b49c40f0",
      x"52b75c8264929c8919a6135bf7e41de7db3b3e4513490cfe43be5d7de4e09991",
      x"430f8a539ffa11d60da882b11c2afdff2cbd88a3c5313d6873c8edf682a028f6",
      x"2bdcf6af8dc3a5603cd52e87441848b1997a2645061a882b0573cfefb435dfaf",
      x"8f521c8dd063b08dcac8636cfb6a8e02d35432f1d5f8a5abee4f6a3ed22cf008",
      x"dc7583bc340a82855c9e2e038d4ac582868eaa1ab9f0abb7b5595807268ddd5e",
      x"2ae721c70142dea772bcf92a1c78fe789e20809f83ead91afad1789932b5f7fb",
      x"a77bc0160ab6d2f24910a3fe6c541de389d760152d0c033f4dcda65e70ed3fb7",
      x"1967d52fadda44c74d42ebf32470454aef7ae0e29f5fa22683e14c533c48a9c0",
      x"ab65d6830317c19cd79a5d6af1faadf38e26e68c1a1591aa0bf1bab14eee4707",
      x"8f2db6aebbf81799f940fbe02d267596198f384f9c86975286e421942eb4cdcd",
      x"d77c1a17d5b09dc8730d924319b41818c8843f4fc30ba74a35c858a3e2b0bfd2",
      x"6ae2942ddc8f9c7420240c63a125599d7c0760c0a7df7440cd7496f85ba41778",
      x"5cb8d92c0db1120ea3ec8212a373e5af203a59674e0e903a3fa9391d71e48bac",
      x"dce31f6b0ce135e4ba3ad8363df1931ebf76bc06f5550757e9c28b55b506b7d3",
      x"1abd7a9c4459b2589d423f4ce32b8621b2dbe05a0f4187db7844cbd0ef06730b",
      x"97c7976e520d2a8e3127129b20e9462732327c57d1f43a8b4248721201cd7a9b",
      x"035baa785106efda89f4bd3a4b583cb2d7e069f6248abc96303dd604115bd755",
      x"0934b1e49d91a021c1b6f382a585eb703e5e76219748d6b71476e66d7c9bb84e",
      x"6871ff6ac75b58cb86f2b760308bfa29696f471e3accab5a5d5581660c33e324",
      x"4774e4be1ce3b9cc39fa1c470ec247f29a3195facedc2e152729f069eaf4bc71",
      x"08b471425fc48918c01d9223c68de34d98444d3f22b4e4ff6a2937389d591361",
      x"d16ac275b774c5312f90bedfb8d661a8a79e98433797f2698a7e9b561a9b731d",
      x"2cd01db713ef3c6e83e1a4c374201c4b46523127bd18ff95f82aa6c60df1d33e",
      x"9edf4fe5bbd510abb36d3d0f2ef066ea7511c55f8e9e745e66432634e477f788",
      x"4d8674048b3c77916bb66486d0c13ea4f18b2a5e17f6b66d08534d85b8965a07",
      x"1f4690fab74d5a72eae09aa318f461a4b69467a9bb3ba9da0433408b26e34ac9",
      x"793a6b1b48e634c6675dd0f642069e97c6bdf5c73067a7de377a78449854cda1",
      x"35cb6c70e5258be27472f0a4c63a4ba4efee9bb0add31ac92765c43b48d84771",
      x"c2f60a668b1c20644860b3b7ca9af1807b0b78c7f667976f11c2cd53e483cc60",
      x"4c027da071db7a19bdf55a73642bce380f50ce3e403d046c081beeeaee87a058",
      x"eb64c0fa63f9db940f761562970e23094d36887ed92620c04e7d91270a4033cc",
      x"9b902d2d699ac6050a800cefefed15ee1a8e396077d50ac626ee502a7e9c6b83",
      x"fcfadc8751ca35c4ff50502f77a17623817f59d4cbd61843078550ea7c4ba0c7",
      x"2c287edc933370bf6837f7ffc4c3556c2ac5606ea65dbd42f82503ac3f1c9942",
      x"d589d67c8ca71c7631d0edc515062cfd79a578ff01ad8ee7e9a6b22ad10d5701",
      x"3facc0a739689ab8b76ab7e663fde0aa13ff76bdb1c74b31a880c251ea317b9d",
      x"64cf81ba662726ede1fb2b6a32144e4c295ae61f3f1d71aed612f381b2f4e202",
      x"be092851eb5a6c659143e180b78c4ef8ff2f5d7057585f8ee129bca2ed4e86b5",
      x"3c964fadf7db4250531ebfbb0ec8974f096fac25bf0cd58330b9c161939e35bc",
      x"4acac941c60ef191e6dca214dcfd75de518bdba2c927eab160592d91ad44bd53",
      x"e3bbfe85e73a67343d286ad26febcdd5924cbde7e85aa43921e16ed1e6f569e3",
      x"823b7f380ae0f5dec7335a15f17c8042e06100b887384370ab339f5993f22c86",
      x"555a719f3daac23503f63b15c00413d462b250ec7a9e8e21e831dcc9f9a4d5d9",
      x"94baeb524a540485052dcd861995132258d6afdd8063af3f9d6b4c404ecebf83"
    ),
    (
      x"2408bc2cbf49af5e51e784784d5f9f1a19f34e9dbd43fd87ce53f2719cc0ac43",
      x"a4516156afe90041515c07bbd15d801bbc1b926d09b3201a92d97d46bd13fcc5",
      x"9f67dc7692eb6bdc11e3646b006bb2af4bb37fd63443ae99a02a6ffe2d5130da",
      x"3e3d06bd50514400900563c86c949db779695fcdd5e8b2d8fd70911c852b4211",
      x"6baea8cf52312c1b45b5b46792b8b7416c45f6a4b9cc2371878b7a3057990645",
      x"e996f59c8b6008c6519dcc085c3a2f4114e0f2499609e92fc58ac3e9f0666e1d",
      x"04fac2c72723d9f2c44829be5940d4594764d5a918eef150ddc5c33eb2081f8e",
      x"a8b8732bcefe775a38642c50f631ecda32b7f4b435b5d02441bf7bcc35a34d05",
      x"df7232d220b54d069f98dc345c9ff15984dc9ebb6942e00bdebac956cc110343",
      x"b013cb8c6112312c923f1a6299daa5469d075e213d5318612189226d0cf86ce7",
      x"96d92cf0583388233a81a6b37d76738a2e09ac62515e38ed94ead38e292c2538",
      x"aaa943ff9721a677035a6fda3fceceb05898e46dd3198635f5ba9967e1c93bc3",
      x"137cc022cd4dbe9b3007a12896a17be4addf956c4497e498548cd196f61fa589",
      x"2e66d1c222f04cdfd33b9d95f06c56e4d712e4a768fce5f1dfb229a540a1a5eb",
      x"187aff605087bdf4225ba56904364f3944d3a7f2c988e9216b456c0ba173fd2e",
      x"eab51d7bd8f2e0871855ed9525447dfb908e57c283ee676d37f5e76afc8cd028",
      x"69f98b6b13f26e82c35a82cc490c5952743707ce2a4930982b280c55af9e6bec",
      x"46c6589ffa6b353fe1ef0341332879b454ef69355e40ca159945726c8704ef9a",
      x"0d12ed9df83aaef469a9ffd210bfbd770260233db18482a57d9b05094b70d421",
      x"1ef3481450cc4c0a32f9a11b11ff28ccbaaaa1e14a893c888ddc96fd6b138443",
      x"84f14f12b466b4f2d86b92b47d7815b8ee4229be167cd8d19ff8aeb75b136e4e",
      x"99c73a647be9c159b80cbfb64147ce4901ced8c8260e5d317c33d1e7970e11ec",
      x"5b3a26c5e41149b6131704be6b91fba857e7f2849e3c0ceec88dc867ca9fe28e",
      x"77bafcbfd4b20b27fa1237ef2f64b44152594276bdd55c0484dce5d4673b965e",
      x"26642e42c096e28f6c44464040a231f6e1ce34ce1cf2c77fc6fa7794336649fa",
      x"dad7fc5d5fddabc9b77f01a40077c07fdb27bc5bb3eb688c3e131752f32515af",
      x"fcaeede016e1f0cf2c0d1908f7d386aac0ff0dd31ad822abe7697dcd78e49795",
      x"447f7f5ef44b822f8d3bedf4c09727459ae584b3ebd02a876edc77ecc4b2653e",
      x"74be56550b6c503971b6aab2eb6039a4b65331eb00964a453962bda554025287",
      x"7f782482cd78300be4a17341ec6bc27cece3195d967a824670a314ecb07098dc",
      x"ea452c260235f681e6ba69deca318ab44829684fc902d01d5bef103f1ab31413",
      x"3d36c7aba4877b1fc254b2bb89eafbc61fa7c7a4308d7470db7d70c55e2ae919",
      x"f9b93868b6dd3a644b710743b950822fb497ad9dacfd8ec0909dd08a70e3bb1e",
      x"1fadedb67970113b49dabc18f2913c3d67b7899764f19a890fb7cfea21b5259c",
      x"c6bada8aec697020a501ea56e1ca9e96e354ca9fb1b40344ba24d523b95a268f",
      x"e494871b6d6bca6c3ba35372c511e429b4ce73a4b42b40b488fba101fe020a3f",
      x"22d0d2f0340c983ea2d481e0a0b8a1257d082eac657b6a1bbe5773fa5aa92664",
      x"a1efa86b2c0478c185e9b2e2448691c90c7bd671c77f93f7eb69048676827515",
      x"0ee272ba6384c50205ce84b5b32fb18f2ce6cb30aad4c37364908e7df10f32c8",
      x"21e05ff36af4c7f3caa34d9db6a1cfc6e98362a79e77b53b7d7c15ffed577c2f",
      x"3d15b5a01d9faae06467fe28f007deec3f4b359f50629bfe061ae6f0c5801673",
      x"96bca8c5f7e09069048b0d76f38916d9ebdd896a0a6f4172fba4321afbc79718",
      x"66f35a2e41eafde3c172d129b3fa9dbbc58645dcbce4f9644a80fae760224dee",
      x"19ba2709263147b671b7ef9a534b667d8b745a436fdaee0d11960b1b1e1c1a3a",
      x"99f6a037030ab06472d216ec680394c266a1fafd3b64442cd2acf0aaf46b1758",
      x"9943c88818e5e09b42449d57e3f8a27beabb67fcdacefe3df305b03535149a0b",
      x"2455cb99f810c0e17f4b98492f964df44a1070379af43d014637cc9ecbbf5fbe",
      x"2066e2f20182273078fdcd6c22f806b3a3d7ba378319060dc004b6d29d58299e",
      x"b4f9e2f8b221a8fd66e2231bb835bbfe22c21b63d3fc29192d14bfb3815605e0",
      x"1bb2e46b1c04339849a24e5b64790dbdd72370193975a358a7db18bbec7fe67d",
      x"c5dc86328bb85c87b929fa0eed250bdd9a599e36629dfeace3ca9460e9c2259f",
      x"a1d13807ce0e781ba07751afc310cc26e302914cea6385fbb1a823d69e4fe445",
      x"9c06639781c5c24eb9545040c9f50bcdef7e245d36ff83c5091e929d3fe2a6a9",
      x"a4f2ee6e892c36688a080eacba413b62a31440c35df7bd81e5812a798acbbd33",
      x"8d3da57c50ebc72a6a3034639103abc062f2b55aefadf1eaafa73746af254d6a",
      x"34d381278ef0a182c1aa94b0258d9f159487e20abbfb47a25ed71637908e11d5",
      x"331802397ef438858d3905d4872e76b2802729d08950c2e4a482c7bd31e314ea",
      x"bbd4b2d8954f79d8a17447fe4538b4ba94ff2ac6121ae538cd351e1c8f63468d",
      x"39ee9767be4bf7caccf9a757ef17c01fd671c2eb7c256a9a21f5edeedbeee8c5",
      x"51447c11f9aae3f198884416bec43ebe08b8bf758d5dc9d0a9d929dc8b4b3cea",
      x"eb45f80436cb3c84cc53dd81e8286fe6d7b6cfc25e16a36b3a02b47dd85d77b1",
      x"70692c011bf2ec243b819cd02e2ba30ebf033328472afe1da8c7a08af4ab16f3",
      x"39c02eaed07fb92b1f70f0d6b7bbc465a61a25802ae4c2bc6e64a1f93cf3f2eb",
      x"69c0f4a660b6c5be4d816ff6c3d165132c9b41924b65442892a6ea15da51accd",
      x"bfd470125e138a400a12dcbe01f5d01fb53bd3028979621de0636aa77c20f184",
      x"35b8bd43f3eca4557ab5ff0b7e7ceb9aeecfae4cc59cf642d2b323b04b9565d4",
      x"4e555567a7e5d1951665b92de09306e9da4cdbe6ed28662bc2790aa8907f13e2",
      x"7c6a5942dd9232cb1c8bcbdedb54c852e5c8470a7fd45c3869fd106f00889390",
      x"0eed0a2796f4d0b598c2eb86043166055984d4b833a5f5ec65d4b9d3f18eb5fd",
      x"f8e5550f39938330a90f28f012ef408a59e090aa67bbc2c55c8f95fd03008d54",
      x"de97384a37a4d0a65d12724db61c29ac7d12ec79a03704df523558d7b582a039",
      x"d6bf10e62f9ca300e6f9aca9aefe45170247fd958dd0b6078b4d25298b656d0b",
      x"dc3e74ef5750221381b2b30a2dc621cfe86a80c9ae542eb5ed6daf2e73e90e5c",
      x"a6631e6b3be8ecbd73d940931d4da0d338ec2b6823f9469f2a130a5d22103834",
      x"3bc7257a3edc0d1ee78fabeb883c84fe9db1cafb2545afbd79ea6c58661e03cf",
      x"d6b405bbe158c75f47c993c9cd4e9f354d6cd10af2fbc14115437abfbde4a08b",
      x"b53e014e9f53e0f940c2819063f065ff7fb7259c83fb0a6c2adef4e85f821e1c",
      x"d6ac65e2850eb00504f6309ed4ac285d09d21d8d0595059a0d020d9dc44dc491",
      x"e2d31e232fb9263c1adc24ab585e41411e054d38976107a4a951199c3e033054",
      x"94c61ef52ced6914c5e355578f05548ab8350c112dccae378b8f56841a025f78",
      x"92047fb2f122e0fac53de03615d6a863876bbcc11ee6ac579cf05576a00609b0",
      x"e05d311fef4e048b95172e5a3f38eb6d728475dbe9a0feb5587f1b4fdd0570b7",
      x"ce78e4b9b3e1289b3e054d4cc0945492b312495add405914c6b44e7cb5fbc0e7",
      x"851b556b057a500e1c82afaa58fa2380c151aa95c354a8b4a052144d352dce7e",
      x"3535490c73dd568c97cf979bbca0e8f5265ad4a21f62330a99fdc9dc2da10aab",
      x"44f6aa6b59483ca921944c23714eb63a8dcc668e37e5e7518c1cab781a8acae1",
      x"a3ffb545af1d1f1187219eb98f69f743c5ead66909e87a0a45b6a3f0868c0ed2",
      x"5f5a29fd8987130fabbd76b70c6f9d40567c1b0a3db538a160043d4fd591b41e",
      x"2a806e995e3b09cb44e47576b01fe152470415bdb0e64c8e8cbd97598e131cbc",
      x"d4f1cb276b3f0c7d1a9c98474a3a652ab87050c53f615c813bd11c1c8b1024f0",
      x"6396a61e6ead2f215688a0fac9a13be438d7a0128af89edf9c5ab70caf95f1eb",
      x"84a5208ce414cc0e79b7f143454154e35c1fb88ee30a7cc442cdbead3c48af0f",
      x"aeb873a60b50c7dcddea9d519c461dff3623dbd8870f98f1ae0cf2e03e5466e1",
      x"c429ee15ad8a0b08ee8e0747b8335910e0b50de018b6850de71cb57da0c34752",
      x"11c257031fa7bc2801d3a860547e8653940e0e4c174c0fe35b11f1cc476a2768",
      x"091aa61aa5b69a863999dae4e9cb26f8dbd4df2386c2e50714fc102feb3fdd95",
      x"e670f23bfd923cbbb026936f689ec8f5c1f079eda5e40a4e9af06a0a49bfef58",
      x"6d534365673d0d9fd279cd955a6ab1126a0551b0df63cdf2f648f31561590db8",
      x"240bdd5607ca128e260ff2ef4434573a750c1cf8d9177ec710bc93d73eb6737f",
      x"f70964532d498009be5846ca78a58aefe369fb5bcfce0a22cc07ba5fe590c9e4",
      x"180b1fac4f11c11925848aab75e2b46ed16963b0591ee428a5681c49679cac74",
      x"4090e2aaf75405952ca9422f6819bc9a0fbd308afdf1ab6584790f6a3e786f8f",
      x"794d5810593c104a72c45051fff64e5dd47f99bf27bb33e7a1f9f5cc9bb07f8e",
      x"e8031dd39c5b474aa147c60bcbac45ebe2b749582e7e02c5bacd888b5ccb7314",
      x"262b4b5e3be527d21aaec62cafea70b4860b79cacbfed926ccc25c07f0f7f835",
      x"e928e94e9be375638faa523f14e226fd8271e62b6e65379c8d54e466d6d931a6",
      x"4b70f8139ef79c2bcce2836e60bbc9319bab555deaa99020245d5f18ec2e602c",
      x"e788a75a911f30759b7778293287663b913cf31dd18e7fdbaa7da943821f1e12",
      x"24ea76bb6c675da61c595e667c12115789fc7fae20169e79ec08e8e46d23b19f",
      x"d62919b7afb5f6168f1686e54b6a61479955fee8c25ebbc248782deeca7bfeb9",
      x"c94bfe86e09610be56333ba6e350b5305fa3fdc1fbd448f5e73fa9fa5131ad58",
      x"b341c25508fc2ec5ab283515f863d92854a57c9be984b33aa19e2eb738574d68",
      x"d9f882edd56d1cc412ed17feeefcefc282bccf80ccac7220aa81e93c9fbac391",
      x"a9567f51624b33f6bf55d7eabcfb2babde8fb6200e4c1af44550da4af47e5d0a",
      x"61c5c7daf1f9125494a2a361d38b4fb84e9e7378d72a2d7f404460a19e901b85",
      x"f003201b2bdc7f72b57c8a36742bf6b256fd1ffd7f950a6150e2d3fa8e503e2f",
      x"94c65b1f5f6848a7bb2392e3bbf24e73ef7d732e8fb2e33eca4b3a1f306b9993",
      x"92aee3302da61c55a29596481dc7e7a310860fc775154d1efe3537f598c58dd4",
      x"cb5f3c6a4d138b3143c1773aabb2c2f6bba6ec2b4ce7cb1e2d0c8581d1eb1f4d",
      x"380fcfd95805a5f09a2702ae2e267db73bcc88b4da11dc5f16f7704bc6b7bfd7",
      x"8bed0b1ec68ab0c17a2a7aa198d5282ccef87797f0e5736c8c06f0c1b8ba2a0b",
      x"c4259a5b72c607c46c7ef0a22e4dd300fbd93560bdb81fef8e3a81d5441cdb0d",
      x"674ff81ea64b393ebbd971d69592bfc0bdecb6ea7eaca9300aaab93e29f9572c",
      x"89aaa41e178016d3424ad7bd625813cf5db95aa614e48b1d08e54557d06ad8e1",
      x"078d162822bb069c6bd073bcd02adf0306f31a019b3661ce9cec3cf7316db524",
      x"65c6b03f343ed6d03b51b8c2cf2da41405cbc830a86b81e45aeee33042729f76",
      x"593dfaba0ac1c1f4f781cb4f0a39f598357dc52b61538d1a8243794ebb06fdac",
      x"9bcef08b0d876ee66732d026b99ebdeb9c9c598c1390ac0fe87b8ef5b16cf864",
      x"1e4c125a06c7251872efcdb8121dfda26c79e6c92f584c8307a7cccd46b8ee22",
      x"23da4b4e3867d1e4f6e9f31951e66c50418d05560731cdca21ff73ab47efe41c",
      x"f43a6abbb80be879ba87f0ac05f606bb8360910fdf6d6e3a8e413da8455edf11",
      x"8f22b4f254f13697ce651ed5742343b71faa707278efae04f840f8b6920c1365",
      x"eeecb900a694075c8cd739ad390b5abf30c36ffba97829f88c15774f7f9d4d82",
      x"2bef765873685394e9458fe9ad445233404bc9d3ef821ed7d4458ed2831440ae",
      x"16e7d212412af8d32ef60d1dace0170e5e9521a62daf98ddcfb8cd3df6b89bdf",
      x"001dbd71ad8ac5648a3f11c20a94a6d96b437e54d61a3bfd3261757d1562c326",
      x"3f47029c56b92ede3d791543db032fe39826286d45c8e9bb1f64bf21ca54c6ee",
      x"d561e27746ddc9fe2b9d2eac215b4052e931aab313f0d59b6bf38c8d2fac38fc",
      x"c108c1e1e455d2f636b1c02679435b0e29d38655142f4cd8fb9a87bce14ac6d9",
      x"889ce823b9152ffefa5d3c7d5d1562ff101ad7563d3d4463f390357ff2e3db10",
      x"3f77d3b1d42bf356fe0f543bd8572defbd1d5f464af43bfeb76abe13e53be4e6",
      x"b7ab7fff5e0c4aebabd9754c42d84000bc2715e460420ce0a218082b17a78b33",
      x"579356f12ee6778f8536075cac8b7e78d11a030f933552125e4990933c59d755",
      x"2e09f71f78a3a4480457c55e0ab167c4da15c8bb5833499eb692409657cb4e5c",
      x"8695c33219627a0912cb9c04f94cd9d0a08e85851b5488dda261aa234de14b98",
      x"e535c54c9470b95944b1eecdbae9b200e24a3181ad58326e4b1d88901c79e091",
      x"60e80b9ca9773488762694e664ce3fa12c72517e7a93ec5162efbf16a1cf4318",
      x"07de61b96fc7e201fd44faf654ba4b0c260d44b64ae865c174fb8f8665180073",
      x"17e81a083705b332027a3b74dfe97f78c26a10cd786f28cc6f25dfb6a6c82564",
      x"f1fd0cf4a04965cd6f2dd59ed68006e3b7bffc9b13f1731cc2e013a80ccbcc46",
      x"a692da903bbc918ff3a7ba46e5a77440b923d1b306c2481a91fd9d9e4928259f",
      x"4919d5c9a24e4729dae4da55c4e01542cd185e18ab012390ba88c3be2a7a4811",
      x"b751c6748183e8ac5019f336c3e04df300d345f17c0cafd094a59200a7afce79",
      x"4ffebdaea22500dc9d037c1883fc4510ec435e799d78ec330fd9db920d6b82c7",
      x"ab02df75ab498f28a385eb24b8800abdc9a40173237d9bee7edf50e2d57cd3f3",
      x"c40ae4b2a7c30c33b621526e40570e3c0d7f6d625010c353a83576ac69fdb65c",
      x"f3e80c2621cf1eb3115442033e5b59517882cbdf34ba700baf447b497450807d",
      x"44d28717f894553df0fb1e9f680c258fca9b51bfa4d971679413a6851969e000",
      x"610270fe0e33cc8870bba166c393024d55b4d6ce17da25f136db51189a48dbac",
      x"db1a42a9df1d4e6eb3fb2ba9f862f5dab20dbab8296cea54fbbafd290a333f33",
      x"771f0eb873194e9a2f19ce651bb84dd937e0b2b2b42e8618844d988a73edffec",
      x"5bdd7f022943486af598f85811433c89a9c3601e16d7cb297cc9a5cd30e37093",
      x"882215223c89d82ba9659a02e70761176d6f4b066c6e4060340b951c8e3f41af",
      x"8b913ed545f0a4e5e50b2c1696ac918ebe07edb09ebdea3c2598ce1999949198",
      x"41266349043c672f4255aabe5df9d7fffc8912a3baaa69861a2bc12e3f6960cf",
      x"270bf2d0afaf474be2289f3092303360a610cb462681d759e285430ac684f217",
      x"d4a33f8b7a17b8f5722ac01a4566054fb3d2f833255c9a6815efc24d2dcef7c1",
      x"b4e6ae94d7257264898478ff5b48c6627460a02ccc8f6e6799f84c2786992858",
      x"4a6e8bfb0e4eeb734423886b42fa8933cc5923a1f626da2bd6b99954601051db",
      x"c2be820bf7306dbd4efc06b562fb91fbe753e1ccbcc6d182d1e2e72a6f6cbd69",
      x"3755cf0a884724b15b206e9ec96fdd28d093359925d657408625334130b196fa",
      x"c86371181c81e4cbfaee915f234206329c6b344f3b0ad9eb2b50ee6969966b9d",
      x"e2d6fd1a4f4e6ae2686a31be35e1134d05994203dd12eeacabb6c16577b122d4",
      x"ff3ebf60b56a7e5d5d03f0297d2c31efb443b374f3f2c6c5e357e73223a208aa",
      x"57da6688ce57088025506f201918e6ccfc5e247db55211919eb4c029becc0991",
      x"423e1f0b8e716c192997b859b6d2c440006cd79a4b64cb3a782436fdffb6f3a5",
      x"b2edeae92a6f80e5f89dd9685f27c4012ac0e7f198c128a430a4fbf70653ce63",
      x"2f61516f5665d72c884ed16ef27fdaf051855e735d612f3b2f482a02d371eb17",
      x"67766749c7473fb30c1d8ba2f5a7e08b4aae5d3e95957b10eaa8f279d1973aa5",
      x"383718abbb3679509f7ebebb3170ffaa61f00900e383f9d231923e6b3c90eb61",
      x"c81215357727b99aef28663a097e9ce0b73b5601303e419ca7cc575caa9c8694",
      x"c1c3a2261527c70fa99bec83aa4d36f74fd21c236eaa43008d2b893346b7b84c",
      x"6293975b54bfd7452fc476e3fe4048826c39f2e4635a7044795a0f4926a3fb75",
      x"b1a354260dbd52f193c716e39d517cccd74e76fbf19168fd9f0c1ccf152ad33c",
      x"ce56adff5b7ec423321de70f3202352338c0eebc61e984255bb470b68b35bfc3",
      x"196c3b652069ed9b5f1bc6d25f98a6d517245203594dd1e97a3f47f6bd2dd383",
      x"a93a11d6975ed716b87383e7791e663ea52f314dd307f10aa19f493d1d7d8804",
      x"66ad842b9e5fa8661966f88b99928854a471484ff84b22e3eb4f2da20ae42dda",
      x"aa8a1fd175c29a285c4b43d5c5f5b940fa7b2b052e3e839233dedf6c6d8c64bc",
      x"dad93cf2773d6ee8a0f92b398f165e65db53e6b6c10aaeb8c933eadb5c7419f9",
      x"04979a42f853ae9e59acb0f3090592398ba593b0d52940ad02219d88acf935c0",
      x"f36b7f8422112cf619f33fd741e43989fffac1e6abc31b0c6ff0488c37c1e958",
      x"33f6973c72a6ad6cb1a57e565bae0a742b692a5423a4ba97e0188462d12bdbb8",
      x"f7dc4ddfef23ab83658520172244248a53e7e029d19a248d0e75a953f4100dd3",
      x"fe1b2d98cd343fe39e0deea91dd9681237cb3726abc1b76a9e0a8349ffc55c9d",
      x"409be010e3d5f233c42588914c62e7baaa813e0b22818f3f8857ff99245d2c07",
      x"6fdcdfe120b5d24fa603791ddc53a6d19922bb3ccec97abfc527c746a2debf61",
      x"ca7c95ef87b11428542d9b8c2faeb131af8f8b23192005da438837d7ba27afc7",
      x"3462ab6f9855a094233cb208a2e07be7ce9d2f2f8f6ddc5fdd843a565faf63e3",
      x"d03c6ab3b5e6f7ff52c011fab2211fa30bb6d9c67f49689b8dba8dc91e0694b6",
      x"c5a3ed333023bf533c43f740c6fa8cff81e66f47703a4756136ea61bd80b605c",
      x"816f4be8f39cde5793ac075455d71bed7f292ea4ecaedc9fb61ee8384551a49d",
      x"4bd7a460b6690c17dbd46c8a12dd7e6d4efbb8bdcabe8a0bef5af2580ebe01a0",
      x"f79bddc4684e5dd02613b289d5d026909bde1fd738e680ea1257fad9e2378da5",
      x"b48a6b1d1694e0e75fb3b6741dbb90fadab7cd41ae33451a0f905adec92d16bc",
      x"688efcdfb7684395741573e702dbe3b4c718fb0495fade5c526e967767aac4a5",
      x"12605949f78389c7383cf87380f6fa85a6884cb2d4409667d4a53b1447a04575",
      x"d6d1a47c610af34e167c1f412778c468c2c93880d63d129d0070930a35be9a60",
      x"9ec837ee5f3d211ee63536f90d0e31c8e5c6e938cf84550de6b2e469cfc0d847",
      x"b32ab7ad0735fb7e4670ab5a78773149b9f0ad837318f6c6c68493f0e20213f6",
      x"81058348545ac1d6eccbe4c2c68328fc20441a1ee663028c09a3342df4104b65",
      x"90c9cfb0b6ab7ae3b4f87919fc0fd6ee9b23623217c4280f2fc8827f6b8261c3",
      x"7ac4ce1fcbb48c1dc89e5e8a7eaac5138d96f57883fe591fbfedc7d1947bd916",
      x"0d10af5c5d432535d1085d8d1a45a63d501049b495b33a23409da70fce70b63f",
      x"f479bd6216a5dd704b05675a7aceb6ee4185e8e22dbd7e062a5fe69139306b97",
      x"fe3edb4faa07202efc88ed613b3c2b35d0e42c6d7634b859439badb7c1fe8148",
      x"9bd7e435699a04a2174778acff94ace390cd4a67d8a5a7802abcdde470fb3ff6",
      x"a79b1a34a0f99213628e6983281ecec7ad305d8b14d79c93bce52afc8f6b1c9e",
      x"c9347f679290a0544e174248b8d06cf5539d914aebca6f40ce06181055267180",
      x"0b1064e2c11270be3290c106642c9242dbf4949ae01990035e6ef6191d6857e6",
      x"23c079d551dad8e833437cca2b6f79e3a566f42858e618a55754d0596cb5c047",
      x"b060b9eb3f15f267c8e4221f97595a9006f388d2d1db07bd0d8a4e0a2ce47580",
      x"628c9e291579b9acb064625192901136ee8e7d52fe9b279aadbc39746df1ff49",
      x"29a489e8eba648f59468ea31e04261606ee748dbf584bd61a561158df903d90a",
      x"c69ec746e41769e7437ad37636a4cba314db458423f753fa681017adee85ae8f",
      x"e146fae85f18cb50f6250c583cfbc29fdfa1ef7f8d23e26a9766b8d8e8399ffd",
      x"06f8fed2d1c7cb16767755eb4fcd0e7e475c301730f846a3ac3a5f92856ce0f6",
      x"1d24559c28169295e748c4cbf053dc4a9cb35faa5e8435d5aac20102b0b2e61f",
      x"4a3bf24f2b2319a3da57a238c26126c92ba90a7c5c344a3a52caa1531aa487b8",
      x"972fb0013f8f6f2c5b4d9308369cb14ecaea9fc208b10e2edffa8d2beac31cd0",
      x"7096f6fbdb525fb6e5dd0369b87003da496aec204e5d3621ecd81b1caee15f18",
      x"a5ea55f00c2e8a0c56c6987f604d5908c8b6377c267ecbbc0a2494d9a44d7636",
      x"4033aba67ca97ec2f063d961519b829f16a5dd5511eeec3ff4262c6b8909f489",
      x"d93ebafee5d5209e80e4d7257bfdc0720dacd9d89d2f4b3361882d75cf2ffb62",
      x"a5bfde6447e78fbea867284812c5449563965806f9d35f911e0ce1de93a85331",
      x"6d1fc95ab0b9b44609f818b04ed1f5fc134ba49094072ce360498d4da0ce052d",
      x"dc48689bd2a5fc9f1af8759a840d615873a42285a45c89dcbd976c6ebff20f33",
      x"36afb2a685fc5e7a695596ec0cc6ebe5437c2cb94b9a037d9c87954dca022fc5",
      x"0c6b4979073d97a08ac848374a042bf8c4cb28f177c058a4e7cc9a2f14adee49",
      x"57ee31bc0e9c7aa60c21a04412dd925807f6774a3533407188ffc47f53b9d116",
      x"72cd34ec42ee35af353d9a6c2881d9bcd71d381c8fce3519d5d9c0cbd718cb46",
      x"8a2e0d40c0914358040e653231bf40c378be496eb1e4e24ad0797dc121e8efd4",
      x"445c6540e9468fed0c68534df955155cdd91e21e5ff2470f62e0a6bbdad8a4cf",
      x"e4447b339418119fea3a8ce92cf5e44bd15d39f197aa5d89f6916baf1a91a6e3",
      x"74694ee04b6bc602553fb9278040f9c1821ed2953296a8689c0ddc7ca5edadf1",
      x"32cd0d0838448f2d874f781d8fb2f197de20b4afe96892faef87dc0f918c3c6d",
      x"1a20a7f8a285c703e88ee9a53d3dc68c29a4e26a7a3b7812f3446bd57ea80659",
      x"ff595f1267c3594454e3d2fe4dd81383c4096913342b0ebb20758bfadc0a94da",
      x"a822a8125d6d9cebbc835abefab3878297f1b92da9aecb59bd38b89ea9fcbd3c",
      x"fafccbc85d6c0e26ef38165f6033aac444c474ff7cbc7cc8134a354bbb591061",
      x"25d35905da58066fa7d79165dfeb263fda97c63687fe89d542a577d371c32e91",
      x"36bb9e43c8382050de8886d6ba6dad432d3b0aa988fd4b353bbb83367c7815c6",
      x"39438a10ea9b095c7cb84ddaf8fd673e14106014a3101eddd9695b339df191df",
      x"1bd8f6c1c9c960fdeefed357b19d06952ba556ff9459444fbbd3a06c6896a4f5",
      x"224fb9cbb31238691ec69d16c228a036b91551ff6bf6d3f683d00f6c1d1cdf46",
      x"c5fd4e3dcc2ad277b5182c431420b2e9fe1d0d6e09906c7b6d7cf358bbfdff1b"
    ),
    (
      x"c668f856a7b9edccd6e93b82f73fc1082affc53e04a2c663ea1b544b87bca625",
      x"2a6ffcbdec7b443325a737ae02ecb6d50547449f15c4cf4c0f33439e5ca93f2d",
      x"ab8068c664f3a56a9dae626d55131d28171b83bde996ee26ea3569c0b9b49ae7",
      x"0cc6c0c312e74c40f603eeaf69ff98bb23238f657082c4c1e6cd8cc640eff9b6",
      x"ef0c0023cb34d5322c530e4b20c85a7029db723f078e0b6e2d0ab97bc0ced6c4",
      x"092b5f666540b8d386f736d1b627d6fc1e4997dc2655b4b655fd90ce28baff8c",
      x"877cfdabe1ef309407cb296d57701d49ac7303dd4e1fe3de3448414c3741400d",
      x"b14492348343d832ef309feab53bb704e6e0cf11edccb2e14ecfddbb2d2b4a53",
      x"3bc0fd442789723e608e64b6f82de33e622d6e966bce12d292b8c8aa3d6e7a58",
      x"aa4cf748b544485ebbaa8a97ca4255f34e98749922bec44ba547f3eb3b8b02c3",
      x"1ddfc8be0c18925dd2f6969aaa536adb9647ecc9fd2ba155fa43b18a42b901bf",
      x"64ea8e8d1f3c4e18b4a0416b375bb227c4c2cb5f31850df397bfc18283887d54",
      x"0559166168fc757513f4ed00e8fd822de1948d9bcd83dcb1affa5cc63b3f8de8",
      x"ec1aee0ab999b062391d1b432f2594ce79680ef207f805bf8a1ddbf33f695c82",
      x"31c51b5ee73dfe620414360a42bab13a192fe31927bc155a307279e52bee6381",
      x"2ef6bf3d12ca191389b8dc9c34d8e99d8589a22f0c9341359b8f0a29a4e04003",
      x"d8bab166e5cc70d0e55b055ea9bca28c381de16c86ac3da7a95b4ece2e1a5f31",
      x"2b2fb33c9b183a78f5269415fab605f19cb05e1c96306acdf4ba423b500dc1f2",
      x"7f6e1e3a715f123b8cab922c51d669d8b24bab6dae4a0e3b7dd3a3e09cb6ed26",
      x"f29ea43b2de2dbc477fe2999e59af6d3e0bc041924191b465ddde439ab7ae11d",
      x"740230756f8018ed55e96a7a065026e25f2c3157bb540ddadd8dc8d782f9bbcf",
      x"5cb9259d7b3a3428063a9511950a0e35c2042a3a3e13a289eedebd1efe15a171",
      x"845fee61606d1b3d12ba0cc720f855281575d08b6a9c7680d50ae62422ffdedc",
      x"1e536b76d848949b5de38ff4360473ac27b29a4a2410ff93e0e47635ef32ba56",
      x"7195804b338c7e1880e5b8361f7f965822551d0b5a11990b3d5deb54e6e29ac8",
      x"7541db98e16bf610a967b22dca3b7e7c35693ef73625d387fc885af9ea5475b0",
      x"37986ca92140b42092693f818551128d8583d62241443330b29de1868655490a",
      x"2b21087aaecf4e4cb74d593159aed2ed30388f60e0dcc74c161eb15759d54bdc",
      x"b7bfe91eb1940dbf7b3e9a1cfb22dda99959702c48e8591d067b47f4149ceb97",
      x"f2779050c554793697bbca1129bf2a2f37a712bcceb8c6bb086b58264a4aa2e0",
      x"c22b1adc9c6af2f6aacf297fe1c410d30bbf387575f2451dc7d772e8e089f938",
      x"79180d7889b85baba9bce5da7676ceb4c712d879d0f3e51353bab975ca161e07",
      x"fbf49a85ebcd66c6af9996839f033381780346f1f66a6f94333a838c19e1c116",
      x"73bcbeec917f00eb6d1a3e01076f764f4921a04bf9729da39a1e82443d48a2f8",
      x"1667245a2c6e767aafda75198da2fd50fff8613af9a1819f71028b51ba9c8325",
      x"7eb6d4953ca3e6ad03c345338cdbec0da52ee3b0222c97cc69de64d32efbd2ff",
      x"2b6e9a9f266bc3b94c31987a9e7a8ff1cc4e56924ea3ee7f758d6de000589c10",
      x"8ac500c6d4e8836531dd29f00363637e117e027d539dde1cee30fcd3349db102",
      x"75e2dabb8ef854be9fb8b623ce2e66e8f134134b75801cca72c19e9444849086",
      x"fb8ca40f0e3a7d3f704fca305b6fee8613127e4a3aea435f30a0bcd73c4b60ad",
      x"c7b9861c9dc45e4608287d4c5e3d1af33978f9d79a69e2842793a21f623f9394",
      x"ae0713fec6ed978bc91d49f4c7514219bec8d881ef97ba0301936c8c57a56976",
      x"2d04e1fa9f31f70c3784b49dab788303e05328721599913d8c65b15bb5b08db1",
      x"6a9f1209842af0f5dec38d9fe17b07ebee8e82c1d3ab7502031783055f381ee0",
      x"e86e030d9bd01d8823176679d0752c6cf13811318885dd192c89db3614f0fcdf",
      x"632a29d4e632a7f7a32a0ae0482204aeb00a57f61e673c231bd52bbbeaf07502",
      x"26dfb00537115062a647d6a46cc4c13b0081743bc71cf65688ce00d6ad0fa804",
      x"a9ba9aca42eae5b58f4eee88e571758f8821c19d9cfaebd1054532dc650dfe59",
      x"4f884798e734c36ae8e4c0692bfa40a7aaec5f51972ddc1ea56050131a1d9e17",
      x"932078e43ba8fd7ed83f9eb91c748ac628020dcb76abd502ea10bffcf13afb3b",
      x"db141d1b61f65a60099091eb0d0878c2e47f86a2dcbb76481ffbc8f2267c2d02",
      x"090f80afbbd5b1c5c21fb027a012e513f5a6db643b1ba57f659d5c36a62cba32",
      x"97be07c702d33ef547ce9a74d3f08d057ede5ac0c58a374ad9bf06b5806af64d",
      x"200849061c515fd9fdcadd01d0d2558e101778dea6890b34f48697df012d4beb",
      x"ef8116b3f5f02e3e25f812c36efa751ed1b01f48085b57be338988e25d080f0d",
      x"c78e7a458adfaee83055056655026285a0b841db147c57e51ddb935895903fdd",
      x"89f719223d99de1b1676c9b14d67a03d14ac5f80a6254c658f92874c85e3e5ba",
      x"748fbdcc43c00a3bab9b0a97d0b62c9531c02e68dad73870802d677aeb33ac89",
      x"d46dd7d39629903748cce83caa803b3746f2a026e8e5e49866577e2f0728eac1",
      x"d58d8bf54c6a5d555ca8b4c62b7ca4650038580a65f58004b55a924783660663",
      x"c0a3c341703bd7a44b8d746a7ac5be4b8758a24afce27f73a733f39b337fff1a",
      x"b8199866befb5269bdc25c238c027b8b44bd1e95588736a478fc9437ab7c50c5",
      x"d47430f9d254e3800758d19012d462b9b84c22558989e73f1e86858dcee9fad8",
      x"ef67f63ce75ad314e7a583e8b4dad4d0aa91bd1e50f9aa22412faa5eac7e1572",
      x"3592aff153bf7888685a3c149d233fddc2cfb9e19b5202e82ff1f3bec312b260",
      x"ad18e5e9bad8d7cd18a4bec37a351e03dbbf791e9056c61922d846cc28d58a3d",
      x"34be8c42956b340dca538f555660c4c8094c256baa45f671cab3610987b9ebd1",
      x"7ee7ef496b67e7866f6d42cd79d4ca185c3ec37111fe256bfa48611ea645fa25",
      x"fef3a1a25596514311eb4fc03106ba8cc1df648772d7986f55630a4a9b79c19a",
      x"760771f270f70fd5322c1c94dd77f796dff4ab7c0f00bde8f96da84233046a2d",
      x"714eff915327bcf0525d17a0c46ef5e79b27f827685cb81463db70f71b90d4c6",
      x"0bbf52756f74bb514457933667e5177209e0156fc33c4b4d1eeb2df9567f94d3",
      x"605cb4910b385cdad45ec9baee4439aea9a1bd35771f8b0307a3370f8efa5dce",
      x"2a8c3e149b271a4a8bfc5b5b3ee3102fb0d9769ee3dee3af0f390d1fb88d7b86",
      x"104ba06dcb955a5368e39f8f86622a28c7835bf26d9c0d5ce20cc56fb8fc5be6",
      x"5b4a11971b1c86e2ae6781a2b0b0c229fd4168d8c9a5c164d03fed763f59f416",
      x"e9ad8d9d287b79d4e88215e97ee13cfb7ddd7dd14c96cf4e716fce86fffdd620",
      x"2148e6d253c73719fbc82c4f673b76e84fd39df9fec3f733f4f8aba664477502",
      x"8c28633037fdbb98554f3047170cb1465e3e0202eb7e22d46ed03a96a3efa034",
      x"80d6199a8fd1fcf3e496fdb2f50995d2a3ed6f673427dc0ce085dddd7541db6d",
      x"e236898129f2360500726b65647d91be444afa13ba16bc6146fffa72e018dfab",
      x"6b5701f9923311a316f2d90a5cf286e6418b6f67683c0a15c685ed01d7f3e815",
      x"e60866683ee7b11544aee8083f8c3b6d6fe8980f93be65c75087fc3e864743c2",
      x"1c2144744a06737199e03a2886143b1981735cb6d52679e55d7536e2b72a2939",
      x"e108a71925c6f0e9b46a43f77c300414dd4ed5901c7138555fa10ae3f11c44e4",
      x"efefb91f645d9a17502b34b5a8d8af0549709c9a81cab4770c7c84a5995d7fb0",
      x"f0e40b35c6ff014941f1b123a70d368bacc5ba536186d3c91f68b18161eb567b",
      x"ef82b9fec2202d354aa4163fd2577d7e9059f427d7d5ac2cc05cc061ce7b775f",
      x"cd47f645df1156d2edf6a47d32a3e99bcd1c926f4d19d03053e4f51eb0e48f4b",
      x"8904d4996ec356b9bdbb2f59bfd13ec90835ee4a7735e279d278efc55518446f",
      x"4453792177276b0e603aa251cf4f87e39fca47da13b5381bf8749f66e9250320",
      x"5eea659cdaab77c1d6e485caf2d60e2a0d8edb767e933a3df33f99fdf3a7e000",
      x"3c23f9158422c8db467ad9a76e0cdf0e9f23ff96f5cc9b72d5392091addc72c5",
      x"904b08d398f0bd8587dfbac69f83e877fa12988a0abf7940a9ba043fa4894b9b",
      x"c2a31e0c834c98e4f021e00e0f8d0392a54af6312bc1a5cf122f5684199750b2",
      x"31c10865f54ea154e5254a5a7671bc0847b4523b82199b8f944ba29ccaca17df",
      x"f80fae5c7f45a067a4c5fe57193ff23f45d6e4c8a0c2fb07fcdd324dba3cc2cf",
      x"501d219061778ffcd0572c8828d0a8cc2a43ac704f18d696278aa8705f32f0a0",
      x"476a503e32caa91c7ae7dbad55e612067fc318f47792dbd1d28501b59d860f70",
      x"062327b56fb56e65722ee7bcd7f2aeb7880cbe247444b9522a40c1f8627af883",
      x"5ff0a92d63b356c1692cf7a7f757cce5297e89f2ba945c67c087355e91f0673a",
      x"f5b42b0cd3c7a728373018abf89318c272ffa4904fa7cc11eccfbec3cb60784e",
      x"0b49f3673b7506223df1e7f4cc75c71d5f0fe2591013f92780b4fbfdd7bab8ab",
      x"2f94e923906217538f9c045566c64f36e7cea71a63fd9a46b3279d80498b2910",
      x"166c367e4c782f766a28ee3fd476e6a095216a0b158dd35083407c99f66cc9bc",
      x"ae96e616cea3536f4a8313d5376e784c7ddff29621fee7f52109297e31b8a629",
      x"c696eb71eb56bf170ab5fea439efb3b83ce3539181c6b7155a22409405ffb9e5",
      x"58df2cb5b9259dba091836611fb48714fb603a9b7e5500f93f3cc644296c1f0d",
      x"45defc029feac1b9bd5cd36be2afcf9bd9d2dbf8d79f55954e4471c02eb67df4",
      x"be36450f3fe9ebb6fe0a15fb00226ad4a17d4b550cff1312d5ee6f4d92786f16",
      x"1e5bf36933753d425906da107ee75d785216af5f9a0cf5788ecc9a91590e4e22",
      x"af3bbb2780908a19454e7160b31f466f33daa044fd5d1d0e19f6e52471512058",
      x"4b177a9ca26bbf1b5b9f3673e2ef94612147aaae7ffbd1b4983486ecc43b1888",
      x"575910dcef1bddc6020126f40e448c1316df59def34a6b0893ddd8457ad3eab3",
      x"eaa21bb7cd30e718aaeff4637f6689d601aab026f3d5fa0cf28d87b49ba03afe",
      x"9cb0bfa04975a270ac0e181ff81838570e8b4503fab518ea1146238299d24592",
      x"13c853d5f675bda29aeed301fb0f7dd0fb019573cd256109c15725591f529ad3",
      x"fdc5c859bf3116cb9df5c0d317c24c2f3cc197ed0e540a736b416cf447f121c3",
      x"c17f7f06199df09021a9bd10158386aef3036c42bf523b0482cfd5f2a49faeb8",
      x"8c6b9b3bee5985823c37f0f2a05ee1cc7fc2233892907881b741e65412ac767e",
      x"821448a3b7699a33b72f8b3db1faeb4e89013262f4d2cc1e646beda422c9cb9a",
      x"b823535a3319bc690820116ae73f7776a4bd3f7d35ec22fa81fef8df0b55ac7f",
      x"36cef5f3576338a04afadfed96973caa8d068a74245ca83d7d9245f1ccaac58a",
      x"c058f1d8490d2dd0dc8e0bdcdf4a4999fae02f912bd6ea994bc6c5db824bd430",
      x"53f53fd5fd3eef49446ccd78a542ea3bbbb69cb21eff823d381b62b4dfec70e6",
      x"01c021a65626fce4a54aeac97157859a3a6bf0d41b9624350e13697cade48b76",
      x"9a50c77da5e9c079b4c6bd9a10aad1e8b6837e0762191c7138d60a713844075a",
      x"01d1639700d619227449fc214b55be1a5c536dd2f1ddaa340d668dbe3427d3e4",
      x"09d174be4182cc640f03df3ca101676e996df387d2e34861d7304fc847a2a067",
      x"2d37a2393715dee4f34838a386fc4e4cd6bc820a33272808f6f9fe2ea4e7f1e0",
      x"cafe026da9c37452c44b9fa31bf162136311b169fc382a60218798803ef1476e",
      x"67abb5e11cbb481633b4b6df383e0209c3db747fd3312511b70e5eda3842898a",
      x"8675a591ec9fb76520676d22709e427e96a03e80520ce675a2ef587970580fe0",
      x"3a458f68c5c47b23a5f9696c24b689b3a870da3e0a9c510311195468f7d0e305",
      x"88529de584269062a6700486e25b3cece098ee8348c7b3ef9d06b585a297a9a4",
      x"d51e8771bc6807ee0eb8bf45b6daa6926981b10913b29365fb87b09236df56f0",
      x"5b4e89327b3bb1d10313994a72eec3e1b6288fa3fefec10a15ccc3e4182b7cad",
      x"ad9ee4e3c628c6eb12582c9a2145e0719490cb94730859f9a52ce976b8b5c600",
      x"aa6076e052c3b8c2a928b4c0b43f340dd03dc367d44d41ecad8ce12ae7a4ad59",
      x"cd940b07bfdc623ca777ddf1c4084f7eef492ba30316552b7b4ca026e80ee730",
      x"4626b4f1cabae43ac4b409824f4ef128e4f4fc6cc1e8b6e7188b889d58040287",
      x"2e860a96020a9c0cfe7af8a4d5dad8e62b7d0c8830a9dce94cba468272dcdec9",
      x"2721ee6f5a19699d7e81c59d1dff5a0a2cbd5b1e56df97073dedff3868ecbe15",
      x"5578c232a3af6be9687c994bcddb3ebb35b1662ae51ae3c3ba0621b9f7adac63",
      x"dbd6a3d53a70e596f132d48872cc2c0bf60db58095bb9a073b7db5f3283179a4",
      x"609798605ec8f8ab3d6d821c1fbfad6ce28d0be4304e696d4d0a3ad74194c32d",
      x"de413d24919ebfd06375e39940416a2ba596496113af898d9e0da9db7bfc3b4e",
      x"31241d405898fa796465b7d06ee0d4e414fbe41d565f3d2ad9f43d8c6a99eaa1",
      x"0d7ff896214db1ea40506e295346d6f8d3d9da611cc1322cc0d82d4eb497d484",
      x"c44bc9a9fa641ed6ab8b16df8fe550ef639d39b61d1ae3d07c3afd6366267edb",
      x"8f9db0601801589d493c9a192f6235268d8e2f0ec92dce012eb5c3a57946f7ff",
      x"c0806a095dc86350e3b20f20e6410ad78929695de6633bd44d372d1ef282a4d0",
      x"6efe127e5044a6ae819c8fd7f426fb187a04669f8eb0e7578d1c98aa7b294bcc",
      x"1d01c0b8c3ff774545f7d6c57050b990638e0462d8d019d0d01e834d0351a161",
      x"aa03ee099c7c9fda328819052851a7b9cab913914b8b09b16730605214924e23",
      x"7738c7cc4b77d654e8a3df2026fe7f691fd75960fda91e0eab4c37a312c5d42e",
      x"702fdb1e1d6c0a0a2994b1cc54e4ea3411bee1f9f97436c9c2bde0a94a719846",
      x"0afe59f63ca781003c2634ffc1cb29589d979c9820c316430643682fd5c95f1b",
      x"5eaff47d92bb11ff9f04a8f9f14ac3f6f53ae29f6de9067b36109d71100c9f9b",
      x"5140f39b312dae13ae2014cf9bb7debe23d18b2332c1533cad20201fadca1cd0",
      x"d507e939c684a90aa462a2148ab02b0e0ee39cce895ddb84289861c36aa416de",
      x"972437f66a97facea2bfca04896adb56cb134f6e6bdd8eeb952d4425c0e9e504",
      x"ff2dd908e7089d549637d6b92bd00986758c555919e2d7523d1a2206b2ea109e",
      x"127fa7e3596db48e67f1d04de4f7c725b7f862110125fc3234ee25f13e1ea50b",
      x"d0972cce0539676290f006bbf59fa2aa707c3b3d1439fc18a0f79effd64e90f9",
      x"31641285766dfc35fe1509cd0f8825d9543db3409dcaf3a2551233a836a8d953",
      x"e3236bd068b626ab6fc64869d6fbe20c63c3fee22d86f1760330f665de52c453",
      x"caded6767f17d82b3c325a1e3ec4b9e2164a57d6e6034f0ccc50063bfc80ada7",
      x"3bc7d1b50b050604603eda3f753704144bb71542faf14a1ef2021cbd5a917c6b",
      x"e0b767a443a15df1d9f8c6c590bb32c72f0fce8ac61b6ab69c0ce184eae571a6",
      x"44eae928bd449137136714a571cfa86a6ea67e31f6968241ba67e1ecb2553cd2",
      x"5c48143fe97794fda9bf89bb4024fe25b02e15960b1df9649cdae7dee28c24d9",
      x"2349a0d1d0d9380671f40d74b0324620692dd19b75862fd509e9fc20feff8faf",
      x"d6a185ca70dc2ddd0b9cfa2ece63e292045f6fc4ea2cfb9cae2ec9663cad2f25",
      x"6194a34bc3e33e9668391be041c31be6af679e0f3e109a36219469e4c9582d8d",
      x"76272723f0febda14a9e68ff41fbda410918b6f7073dba819a720915e7acb1e1",
      x"94ef58c39dd73762a223058b41bdcf3c689311ce5b4558bc76c47930575ad568",
      x"94f6eed1f83826f49785a90d6dd385c9d324553b03b74068f52e64d79802662f",
      x"0a1fe739cdbd2da7bfa7244e1e9462ccdfc554fe943bbe5c3627559859ecb311",
      x"ff0718d3ca8c1a5c31dd1b82babf6ee6e15209b56ba08d4c1895fa3e87064a75",
      x"56f68e98905af5286a9cb3480746d9c979c629f24d4164d2816a98d3e59f3da8",
      x"af92f62903d46f989b79b7ed44f7e41c9ca6e5c90b8c2ec8c3c2eb4d833c3b9a",
      x"c235f87044d038ce1e2f6ab78769463c85d28a98aa7d7d78553e3e42038ca7b1",
      x"6d725cc83ba45c0ed48066fc3dd8dc45f22d7b5f80449f2f822175d0d9283402",
      x"f73a25405bb55793ab1997f1f3a151e6a2aaaeef0e28e7207caeaa3ca1039798",
      x"8555ecbcc36893f68aca5d87591157a34d32f0c072698a7d0da645fa3bd52f09",
      x"cb7f681c17310955c0b87f1547dbfc24282128eed99e21603d2c3ce4d06e614b",
      x"1d3a6b9e41250f5087f732f4a20f61fd7f707164872f26740dd4a8eaba37fa0d",
      x"607650c3b0e1b851fe5b43f22cbde8110ef666ac6f3b2ede9ab2d7abf27bc961",
      x"231056e42ae8001c0c99a77af8f27c369b7791f3c5bfe456e8d74eacb62e1c3d",
      x"3f57090afea751c5af0762126e8e9e641e73c87d4c1d1426d98a1a55db428e1e",
      x"03c74b122cea9c23f378b7334ccb97f852f20d4e9cb611d029c72f5e3f1f2749",
      x"c30fe6814430682540196111ef9efe97b90985d889f3c90e8b4f568c864d5381",
      x"852052088a26931a42d603a10696cb89e44ea31cc219065f8da61645019cbd36",
      x"4b5ec9b2f97eb926ec55069b8deb258ea075a5b43eef7f134f030763f9fad83e",
      x"00189d271084b4279dfd89e946d2da2d8a5a963c7ce1c45f016c13d7902dbb76",
      x"57fbf060aa1e355ef44950e36c588f31fe18e66c7c3637ec151409269dff08ec",
      x"9b718e10091efce0cc573969cb6f1d3684c21279bff7dd1c82e5c5d5d7018912",
      x"f53a84537c8d65a12235a817c680664aed47b99f32ca2b584c55442b9ea7970c",
      x"cb1183d25e0fd7d7572f6be21fd9909fec8f0155801edf9e6970d511633a3a67",
      x"38af6d3494786d57896b503234b3995851a59fa316a6ee93159edd5b22a85082",
      x"27ac8300443db9344c75bcc8f3bfc5dc525bac1843547867f121efb190eebbba",
      x"f80394a2fa3ade345e56d81fbe0776b97b3245f2a0861178cef06ced2f5fd98c",
      x"bf1bf870ead3f0073a16cd3e27ae941ef920422cd4f43c2504605fe5818be34c",
      x"e94d7132748951cc70de672c0a5334b4b929ac623ad8829bacb1a143b049f860",
      x"c29495b5929473df52168959ef2642861ac9f3ba6edb1cf30c9a474a1a559289",
      x"47809b21c569d2100ff583fc0545c71d02fa71128197824e3767c4eb496d16bf",
      x"5f91a18d45d552b3ec63d56995d1d67ee3517e1392770ea8ed752ac3389eab82",
      x"c256db2072d44de496b2c5f94644d8ad92699c7a3becd85931c6b2db8daf7ffe",
      x"19c050cdb0724bca1592db9b53835d41088e2d8f393ece3106787ae732103b54",
      x"da5bf3e3a105e56f61670d540b836ad8ecf61643dd6f48d9aa9c4dbb8c019cda",
      x"c8a7fb8fc9733fa7f4d8882449f57932ba46a1588c7779e6d614d99c23ab6081",
      x"cd27553aa7a5d6260edd080620339b113a5806d86258dbbfc3b66a1004858ff5",
      x"bc496be927d505d841f3ada11a3e561ac991da8f8bd4d45086465eecb719ee70",
      x"24ab64bf70e187225c37a926822e505e22d54993d90038ed801146944582834d",
      x"bd0e3d5933c1a3e92ecb2e88309378031e597482f2233c8695bf1a10b13ebc45",
      x"7ffb85c6307023fa9c67c7bcbdf87c42d8eaede461a364eddb437020fd4f29f6",
      x"6957ec5f453672d0fce6bbeda450977ee4001c6b4949fa6cf7fafa7c4c81d72d",
      x"ddac9ec406112ddca1329b23e12f4db46470bb86d7c7f144e4e919b6a39d3fac",
      x"c6999ca1ae2afdf789158ebb6b94d0ab4b3989355f0c379c34438aa82347b8a2",
      x"49f576f565088b85c76e5894d150bf9199deefff0af013e5b9086e6dc0382747",
      x"c9b179a2ade285844e1c6edeb054d3162803f82225f34286804069a4c27289cc",
      x"1475c4db2ed9ffa503255306fbc3e82f45027b75e112428d3d9c7fe33f1998ef",
      x"927eb96df5154add4e6b90cc18f0e5de8f83d2fc2f3786a0f6ae0e22b1213824",
      x"d7ce58f0a9617d7800962603c216af59d54a39689b9d7831d1346f07162b0d5c",
      x"bcb88129dd89d47845b4a27578267836416cbaf82a28d5f1eabd011ad1a0bfd8",
      x"29467fdcdfc78f4138e55c4d6340030ccdf95d6bd02078dffb0a9ec872c99046",
      x"9317a245388f054dd7e337f73de0c8ff7ad7d892fd0e22ea852fb6a6742deba2",
      x"ea0ba1df2d4689fa0022428b23b2b9d612a5cb36fe41b951fbf1616eee2ae5fb",
      x"9544a1597ae280a391457252e833c6c483eea3d00f5c666e7455c48e46004131",
      x"f8d66603e49afdbd3eab17bf3ea6f614200e7995ff38fa3becc5369e73adac57",
      x"702aac3c839d7e029ed2f253db722ea9cbd85228f502ead40cd7774b43d8eb8a",
      x"9aead3f98a3089ea912bb70bdf64faac2f2beb01916bae92dd0b25294c1879b4",
      x"ed234b7abfaef3723c0bfcacd0615e0316f37ce32cf3a5c38f57e6a822b225b5",
      x"9998f98cb18561a2154f1fd0e3bc7931f6919d14e7c9e8243647388d765cbc7d",
      x"d8425dffc9a5b3579df663b2ea7ae18b7b0125a9ff750b76d56370d521a83ff7",
      x"afa0800390168e161cc2c39aba98389a50c9348b683b69072b7dcb6746e512ae",
      x"732cf7c6b27abdfd2c6b138edf94c5f2e90beec611486d2d835fe477131718fb",
      x"2b30ed8c9e716bd5def44c087a30b0127672a367421fb6375eba75f8756cbc74",
      x"307057ee65979184c7351c97c5203e15bc402a160e3ebeb166cafb6ab8c58755",
      x"aa2164673632905ba56bc28cb1ee0ac9c3286a7051df35624af9bf2edf92c45b",
      x"3341aa15748a6485e184a26429bf2f3d81aa9e40271eab49dfb77ccfc2bc218f",
      x"262731f27ebcdc33baae238be2868c7477acd9ba5c5ca542e1d41cb616cf1ad2",
      x"2d7a27101ee3e765e50db14de86b0ebe208e11ef1c34b82e8a87cabd318271ee",
      x"cd3701982afbbee77b5ec45b497270f2e6b76513ea14b9f2aae6e19801ed9007",
      x"e402951431b51dc694d519ff462f993d539c0fd31dc3ed08589855ff73e42fc0",
      x"c9e4a60a17b7e8961ccf47f7f567b61a7132ba59a050e65782812a3327b92bbd",
      x"27c6550c4bcf6c04f067b6721cd12cd6725ee2cafc053414a07eed23ca714acc",
      x"44f8ef559a94c85ef84875f548ae5ab93b07ac4e1b91347bc5e37b17c912da65",
      x"7b990a27bcac7bee64b76dc03022ad773521e202adc3906a5e0f06d59c61a6fb",
      x"6ed2d6ea3620cfb3ee80f36f1494630ef478e45aabb23e34c3544bd4ded3e552",
      x"1a07d55225c388325cd67110bde945a5f41df345362827f6dc7474c0f5d1e084",
      x"6e7aded2f8f0aeb72bd8e26e48ec65b40e9d7e2e6965b7710cc4d29ddb60a1d6",
      x"882838b53e59ad3188cb5d834021d2dffda23f8626bf34c8905477b178e54228",
      x"b11df438e73225e1398b66611ab87c4a200cf3e32d80da729e5cf48fd05eca8d",
      x"cb63864dbdfd34bd3a35052b0c357c4aa80558f256a98df1d891fc4f2fdaa868"
    ),
    (
      x"f356d845a33419a0fc3c4f8d09dc73201f3886696df6d432d576710b1b8f839f",
      x"675ff4f76e1e5160fd7fba63160d9e3dca406a3297f5301161172272e8c8af7f",
      x"d40fc32bf38cab5f139de60c65969d50cd9e4c9acba5fb478e16dcee148a7630",
      x"ab35ea919775963f0b8477ff26e9cbe912268f0d3b49524dd78e345d7edf6437",
      x"fcf0051996e3f057d747810cdf39d785f889ed1bc52c2e3411765a3414d22f57",
      x"6c7e46bc9dc78cf1a5804ea7c87ebf7a25d661812ef8777f892f7f5478b39a23",
      x"9b8a7095a0cbd5b661ae5eba698ac6535cec118c54e9b4dfb7aecd65a83b0096",
      x"10fd39d56e9203cf961790272d289b15a2319ba439b33c080946632a9e7ab9cb",
      x"055ef51e3af60c4f97c4c5868b9c623d5c9a61bd10177c2a900a745f39b32cbf",
      x"0ddeaaba2babc99221b08a765735cfb8c6ffa19c9acf748e07a32405839b6e3c",
      x"a750d8819103c334d734e2866aca5d56ebdc1a3dee92d89e496cd6bca0690da7",
      x"e62d43e9bffedd826e0548f1c2a96cc1347934768863aa6566e7baeaa17db655",
      x"8d91df70b93638319e6334d7b2eac3117fa88c0e6b27522ccc288a1b4a3590f8",
      x"b53a79e6f4e2b45aa5730769d1e64d7faea3a22dfa062cf8a73ed3ead1d72105",
      x"5893f46d8f23d5c94447db0b7cfaeb6217e5c29fc35cf5aa96af46d0051094b6",
      x"fff2e69accd6b28bf019072e4ff9f1a6d040ea8e7b788eb528eb595fe169ea11",
      x"48d2c378f3092bb65ba0d77d13f2ede48fbeddd4c67ed5ca5c7057c6c20e3120",
      x"844fcdbb87edbc22888b3c15ae64f040dbf919319327e5e227210652711abc98",
      x"3c66d2632ad99ce88f7f0a8b441e4ee7d83f677546ca9ce28e6753b88334ba1d",
      x"3559cc15a720693ebf129879a3bd07bd805764a54ff31d86c139191bee9e190b",
      x"1ff55a68be1081e14c6fe9a186b55b8ffde83ac816ca75bebe38e43dc6204619",
      x"7c02871dd4e385c3be3eedc867fd96bc5d38068926f8c49fe034a7e446b48a75",
      x"5ecb52e984d7faa8f87a7adc9a1644aa1ff56edd31027f4e1e612df4bc4c0563",
      x"ea3a2dd4f865606128ab93bb6842cffd25d57b401e8bf29e243931c658c548e2",
      x"848d43f91ad40871979fb055134c0c0ecc4b7863d21a51745fb2c623dff5bec2",
      x"87a961dd9ff781bf204562da859a13cca25cadaa83cbb29a9445be1a08b33f6a",
      x"4d9d051e144310f6087972ff7370af053683ecc05554e2a42809e59a4f15f8b6",
      x"730012c490ecb83dc87555110cfee49c79c707272254408b2724982a696bd36e",
      x"2c5da530d7efe1de949d0a572ee7ec500d94d5206896c0d0a1a455345094de03",
      x"09a8be34ff799ebfcbb31eadd56963b9083eb8f8bc4e3533ae23f93bca4eeae6",
      x"922b1f8167877e3e6fadfe0a82efd7733a5ae416af477a3716225d6883c2fffc",
      x"9b924f87c913188f74ce31f5fd9c77154c59d746c5ae04253378c9512e884374",
      x"98e1c0e163ca6581a76ffa1523d4a8b5b8a1c54e6a2906997025f4e7aa38a356",
      x"b947bda6d0ca4fa107e9241909bb2b4934444800eee861f8475bb9d078569939",
      x"c353508fc056a22998294a0cfac9e7b913ffcbb965d2c5fbf604f8263705e806",
      x"556e8242bf348f3d325e8f5b8bf631d7766ebb4780e95ae1f06a298bc67848bb",
      x"c3a8e4100e12383ad8b16408f714988d9f33bee4961fd1de2808980c6705f131",
      x"1d743e20f26a559eb89ec42f5f54fed3bf89beeb9b85ab3156fbeffba2812e1b",
      x"8bdad85ccac5371fe5bac12a0b98a8c8bc2345d34042c0c59dbb427997409c81",
      x"d1b383bae4ef4d4b440cba136b22767f0b0ea20ccd90242b297968a827a8c757",
      x"91bf0444936fbdcee50ff4164e40b3a63af99c4a2462636c23c3f66887d0b767",
      x"a617a20de16752ff989ab6c8c22d3336bcccda5f90f7e7c7b76bb83a507d585b",
      x"c3c0fb03dee58eaa0e20672a44a0bc2c67bb809e1b29345e334c328908d28de1",
      x"968f803bb06b71dd2d5d7c6fa578fdc2cd472d570ed00617ceb1959b1869672a",
      x"84d7deb80569805896120e14a789de726b5752406272b74a733eb6899cbb6889",
      x"224529bfd50929778b00a954c53dc5b9a8f43bf3ea0d8a88fe6421495aaaf871",
      x"4396ffd49f701ee30f11018b418095c5b3ab4842b033c04c54c5476f130926b2",
      x"033c69eea2185a2fa8d59325c267add5e97488454f325fdd25c272563b82944b",
      x"a29f65d891428077cf0b245dfac2f2c67cc88c3e28cc789e10a8307451963ce0",
      x"23bc23e32299b9b2fa380935669704da1cc1902cf8711057c6f944b5e38e9a6d",
      x"069446ef7abbc0fe046e6fabdfea5f3d8bbb1663a21f00e1215f5841ad97de57",
      x"5f1ade6dacb502177a0753b9c8e9e27b1cd4304d490b8ba29b032b55fd96e2ec",
      x"efdad3c6a9cacee5c47576274ab6f8cf73bb47dc110798bae3df7e5b14533c46",
      x"71100c6b040541567987e8d83cce2e8f7b27ea82d58aa995c1c0903777797d45",
      x"21e7eed29f05e712f787bcf5c53d7ec71ce61446c3ccf6225562957ad159c36e",
      x"725cd3daa8071aba8cd59104b0f72d68799186b9968f0c1907c3d93a777e0ddd",
      x"5a3f1ba4d87cca1dc5678d0586d36da5fba27349800fc3fcab306cb905cd203e",
      x"78ef28fff18e4c146d8d9d9ea54b91a16ba84bd589966fe0dbcf08fa5af67c61",
      x"ca575099b06ddc94606ed021405e7f9d46e9686e5ffbc69b76e8214d8add363c",
      x"9c8512310f8156119a68f60132c6d1db108f4deb6ad55755fffcc47a0d073606",
      x"68e2f03dfa50c648da6d6fc7f8e347fcec32766db3c5f33e0195c22f466d1ba4",
      x"86c460b7e96e158522a23b19c95fc357e0633dbf054284775f8796b8745a1916",
      x"bd4961d81bc087d4f22ed95a60bec81bc43c5f63c23001fa7e4d505fa36e6b8e",
      x"a55a49421c32728d08df29b55971471ba60c5bb687d213b53a6f77537ec6d37d",
      x"83b508164bea44cf6923fc9cdb4fc1752071bcbe59c5de84a52e3e931a59558b",
      x"eb98bfedc60402059000024a51187d5c2c3a1d5c700f6852596d875850332e6c",
      x"df8be8647ef2211a5b2c97534aa2f1006320664c793ec56d3648d90f7f3d64e0",
      x"06e02ba85e974a4403e9f12f455ebff0de33c70ae5acce532dbe66bd2a1c76c5",
      x"6a12788f11c45f57bd4b30c42bf578af782588908a24a33fb0088fee91183acc",
      x"4835733ccfc922479d9c2d51eef003270150aa2798f429a20d50f763a673514a",
      x"a944480c6542ca44485fefda50161f6e06b0011554ef121e147273dcb45a8302",
      x"8b024cc9469f3aa1109e2572b6c243aeaeae6efe0b2c190a9277f537f51f1ad6",
      x"1e115fc77c8070831786f3f39fb078f4839a23fee30146a8132da75920c131c9",
      x"ffde0499e16dcfd434501b7013b9d84e8bf3faa353d2fd2cb9772bbf2728cf05",
      x"ccf09cc55c550885a811b63d3d6ad095cf7a624805c115dcdbe39b90194b4bda",
      x"ee78b2fd990a4c93490f844b8651d08ebfb8f4492f38ecd34bfc8c9110816d6b",
      x"817658f7fd05676d189a17db74910204f7014f78b0f1e6323fa3947a3630c9fb",
      x"0ea6ec7652b8670041ddf0c84a3b38a98812399433bb7d033009628e8afdf447",
      x"37e00215875ef65e36c81af0dd090a911535785d5103f1997c50ef8a8985d781",
      x"b28d8f8e5bfb626f17576e3835091ac0deea0e05cb7d7d902c8de729694c4f36",
      x"4b8fb6356d9636095da0aa697ea4d75a6de32f12d5e4d0268a1d34be70445993",
      x"3f1b707e0a5654ae19ea7713816b726d9a52d30beb645e0731dda731839687b6",
      x"52543ba637fb8e2ef9c56858ad833120187648788f3a036a9cd11c6ad6fcbc3f",
      x"95e22dd6aadb73e77391dca6a52a3a571942c99413e29068196d4a8403b33e85",
      x"58ccf63703665cd8bad37af5f82e956009ecbccf16bf63b26597961714035d99",
      x"5b6fa7d9b714274c36392d1aa8fe29e197bb53511c8f618bcf8cb87279e0d2dc",
      x"a693105a35340afdc92b96d5a1e72ef4073a868b66cdbb7889e861705d8c264f",
      x"7bc87942a3e8a32d26119c205fe43957bf6cba2502e6fe0bb44f58b06439a5dd",
      x"5e74515a65a6f71eaf112aaa2ee1ff27c75ef23bef4f7b9bb9be424b11a67769",
      x"42947e5e2017d96dc3792ce18b659940129b50f9d4ef48c4c9af2575dcde71d7",
      x"31603f8d9ef33fe9a8da885b872cd01230475c65189802b28c35e1bc446df7f6",
      x"d3a036d7d0f1caf444ee65e18711b77c9dadf383150a3c2286adf003ae5ec798",
      x"781d26a01d82f1dfb20def93b9d2de84b9582e4afb349b2c55c90a726e7cf30d",
      x"ddfefa2cb3615cf463698665a2964f04204e27184cff68596e3985afca1fe5f6",
      x"180bc7b1ba26540ab93d05099e093206534d646e2206e8036a301ef926eb0b61",
      x"0bc30f133a0aaf471c411e05cc386c8df1ae1e2db745573e925f7b6c594161bd",
      x"7dd487e3435d3f8516ac07814686e1dde929957ba71e2c50a5ff438d62c67073",
      x"332bd6a362852fe730a9771c85da5ff01bfcb11c0d99a10769c7da26715cf3dd",
      x"62bf314b7e65377d1173267754fdb3647aef635beb78f4b1dd7d1f446a86fde4",
      x"8ac4563c332b9220c3721d9bec30fb4b10b79e965682a81c332b63e9200640b4",
      x"3aced422e0299bbddac8b7459ba1bd78fba4e5d7eb73ca5c812b535100159c55",
      x"f4933feaf1f2962a636f1069016e5173e2da7ce0e51246dbbc2825897da933a8",
      x"350c6fc562d2b3f11ef00675525162779e8a96a1558ad697bf5a07255451aa58",
      x"ec001874f66636f2694d99f3c17f7b30ac7c87b363922569b112647e213aac2c",
      x"2393aa6839674078dd42b722501e4070613a1e6475f36487cb2dc5de91cf96e4",
      x"df6374152761256e57250b7ed0b8c39f70a42dc00236473de0c06678da27d575",
      x"56f6b69a94ae79dc14f66c4735ee1d3c3d2f6a5f77399bbc0d2bc04dfd1a60bb",
      x"5323d4531835d0a27e5c0cb52843f75d170ab3dc287ced8834d748b05a3f3f0f",
      x"7b4411a13ae202f6afd468cc3b064559c4031864ba89542a65d4d1eb3ef14fb8",
      x"2b92dbee8669d23eb94999c3c272580f71c4fb72cbf4cbe02013cceb058b7a8d",
      x"e53f4bb8d05e58cbc39bebe7db3086504cd706fd3b2338484fcf76ba5cabedbe",
      x"8ec5712f74a2c3944b9f39c98e70e1606258555f52a4292ab640d13d04ad2ec6",
      x"8f6f8bf292be80e5b76c5a12e58fe94db36133caed7982ad83494b4fbb081c34",
      x"21f371eea5069f31d958db29b37e98847266582c93cd4083c57ed32abe7c37e7",
      x"c57d740dcf7045a15126ca846fdb406d263455990df00512182c464bf28e9e16",
      x"eb9cc8eca784aff160ca163e944eb5eb0d4d80e08770f18001e7e9e5e67244b2",
      x"1a99cb5a2d228864e8cd10e6a066d302c5e54c5918b11d85e4511e77cf8de247",
      x"33a5905e5749700d16f265372feb936626f05cc1561f59d40d6846db5261c164",
      x"9e607ca56293aac7234133ec4279944d6cc9ff75309f32a61e0eb3374b0d2f1f",
      x"17a9216d62246f5bf2619be4d5a0e473d5284415da93d8e1854127a7bce80836",
      x"3e25e4bd3f47028ac1e6c2286d765639f007c82c95b783ed5d1d085b0e124861",
      x"c2b61a22304538c04bf586bbc1a103542a10ca32be797911a9bba295063fcc4f",
      x"b7d6325eaa5b0bc6bd70227796e2d369025121f2b0861733d47b3e4d6e3e910c",
      x"dabfa623549226cc647e30cec30f68d13112d6d84127a5316b5468c149572913",
      x"82e0487e5f923671c13016c41c1e45ccc5a239b7b65299d4cc35dcd4e4fd3a56",
      x"999926c8e4ef4194e8f5f95342c2e6258ff534af4bfa7ed1a5c28ca04580c9cc",
      x"8c573b06ee18f582e452ca5f5bb68dd24e907cc8a6364cb3f048d15e30555c91",
      x"0f328212dd8a908f6198103c008070e35b6ef7680cec06efc5441105ac6cdb0a",
      x"94b2c98576d5b98c28a3975a61027a5cd467b4439631ce23e132d3984e6ba93c",
      x"3246f06f7ac5cd4e555f3205cdbb95aa67fc322cb87a4656959d1deb061005bc",
      x"cdfe87e0583aa4ca11ae13de79f7f1e6d18382f2644ac35a0cc3f78e4a307cf0",
      x"0a4d6b2add6c9ee6488f822693e61b5a2dc23ad99040b4633d2bcff6dfb3a80e",
      x"912dfeb58838c83456a5a445d60a6f266e5fc8b18b013b986a193b2838c772dc",
      x"d3dcf1e23d7783923674a2b87ac0e46e04741ad91935d040dad2a1d0a6228c20",
      x"037c8bd09e54d71039c427e02df516fcce67a6137c9ddb1e854c7d063f87ff86",
      x"8d3b98e23959135b196196b079f96640ee66b39eccd1e6af50df09cf4b59af40",
      x"2aa978ec76a9d0f95d0b9dd7a18021361c7654da841cb4bebe80ef704ab655b4",
      x"a9e152031f4bbd577ccd486af530800a11bfe2b9876d35b039c109423e7d3939",
      x"b64a9383ec60fe4250603f87733863fa7bbc48929812351bb34f2d70ec4a36b0",
      x"290f95c5893ec29886ddf194c559651edbae01cc8cfc054a38d6dc93440e96b3",
      x"ea53eb764de995d92ec2faa6527a30bd8fcb846ef9c2f8e0a932b49b62e4f2c4",
      x"89cf3dac6664e90c51a60f597b04500ce3a6e64c35daf02320557c1b900fe567",
      x"7396ea25cb2201b23d4568a48a1fab886d0839a931c988398fdc44accab6962d",
      x"473db5ca6f13b9aa504b7c445f69d3f87e624f1cfd2d18075898f043bcf532a3",
      x"7b9e39b178a02888ae7f504526cd43a9cf927010ddfbe3864c291e118a67170a",
      x"9159768b936a5f49e320d3a5a03f46f1b978f28ccdb51d05daf7567bd4e427ae",
      x"177d767c3dcb8e82d3729b3aadae2b4508d8dbde3df5aa2941182c0cd9ca5ab3",
      x"e083e38873d0810a4ffca3d7b1cb098a49ff07bf294cca3dbd3d7c1ca5033e48",
      x"b62ca55caf9d1253d221fda77d288b92f8b39ac596c8ddf49c2c8b39ddbd57bf",
      x"efb03abfdb089b963437c43d2dd01eb4e7ced253010750b812a21f5cde9125fd",
      x"c298d581898b043dbec0bc267e6ccde903e81a525661964ff66e757199ce750f",
      x"46638e5ac185d2a85fc1d2823f91befe9f403f93197041b5a528626675e9e7a3",
      x"7c1c0579fedc83c1845933a375811852e01d3768b083a00ed61477e6349bc600",
      x"8881db5d9e400166413c1131d8a11bd617b12f39053d01f2b2600f7c9bfc8966",
      x"1e73cc2ee3e14e40937f6b8819c85fbdddd58c322ad70eb1aa65c9e526cfc563",
      x"3a1c59ff32e8e8b4da94970c338d20894be2e57ed24053004d9b5c82d8543743",
      x"47e4532a227058825b089a70fe53c0330990a31701201d2f2b79af743bb96a43",
      x"da87da3debdb8f05e44e6fdddcba33a1725a94e686d4244bb493509a4ce3482f",
      x"b95bf80639137aaeb0831f2bffa657de82393ce0aebf267c9eb60fa82afa60d9",
      x"17e7dfb04ccfd2e51b017a0912bec9494a9c860a1fc3927fd4d169aec819e374",
      x"d98d923e7a8270282fb1794751c3f8b6a5225b55e55eaad0a7e49265fd2dd3eb",
      x"69a2c46a89e5febfe16d4e2d708169fb6a210dbd0011f31e3d3a5896b792ce53",
      x"18053cb0ee8e1367acd7fe85d7df4108b662d01ab7e82907078aa29bb602d8fb",
      x"5ab118e433d47ebe85fa9e1799c8287a248f6b96089c97ec029978084cdd3f07",
      x"ec7e041d373a40bcb1bd6f55a0ffeb19031e3a5868dcc6485f43faa6ffc8d525",
      x"03dd8683cb01233f331509952d7ab761db2591fe4d1c5edd01d6eb16192a3bf5",
      x"ab296b3f6410070d15f5783c2efc9660427a7658162002381bae9f58bf3cba46",
      x"2b8599376951d343b20810501d8b2587ef9241e6a45fe3d8b54491451ef87fa8",
      x"1e9f20c0c070621608e4b7b77bd78bae010aaed5d91a6744bb5379c92dd9b120",
      x"cffdde0c60ecdb84c04e2f561b832ecf6066cfac1b412eda5ab8a6eb120aaf89",
      x"d14f7449d9234890bf070f1941504c8db118ffff103b3b10fc21d878521a5415",
      x"fff66126ad84507713d98c11cbdef0526b199e9f52096525023572a5212ab383",
      x"854e761b7e0cf04069dc813aac34cfd72156a03a0f26e717fb7049b19f1b57ec",
      x"b8e4ff76d85479120b63cf59ba31889287431724600ba670f7fd803be2e39fce",
      x"e165be1411353d4de07ec76ad6f465cfe4155de7e0bfe8d80edec0e17a159e0a",
      x"af93f95da9f854f89d5d3cfb55700ad828d34d21c80d4c8c5abb267aee2e51bc",
      x"49eb930bc1030ae40a292234f5c302e055738be88dd0d5b8a922a31e65704d81",
      x"c9ad8b7e80aaa634472a8eae0a86f4b55670f6ee74db46fa47be789db2022ac9",
      x"4f2784026457672186682c4f10ffa6d425993e5eeb3c1fde4090f62610311520",
      x"2d542a5d6de0a991febae21a987ca768e0366c9b593736531ea2def71b44e279",
      x"8c0dccc61f88476293a8eee8fbee3aa902243d047372731f9aa0df8272b81e0f",
      x"f660aa083b6dc38bd15effd13ba64e7866ead2ac8c9e7f229e6a86e0b49c6f4a",
      x"0a79a3fb2a71907e332d6a98e63735bc8e4bc7ed6bd4918cdb5e46d301c70ab9",
      x"1c98bd7c056844caaf6519a27d1ed71f2cfe1b7fd5e179293abf22a68c904d52",
      x"374f65912344edf066533414c573a008ca0374bb3df21d8222df0a1f65143fa3",
      x"bd7f5454fc0cf66f8cf1c0717a22a96e7e402560dc8555944519b804291c0769",
      x"d11ac4fc0a4a171fae151ac7f2ad3c3064659cfff7c8dcbdff0baaea4139c3f6",
      x"65a9489a98201c3d0b8b2db6064a76ad51d8045f6c2adf5478bf38adef5e6ca1",
      x"3356c6b821e15eeb0b541d4cdec16d0a7db6cfbf27479be5b9276f06f0a6f725",
      x"428600fb65376a1e75a283c21ce786e993579f848b8594f60fda7d9b0bac005f",
      x"433d90b347e23edfdad633ddde32081886ef8519c6ecf91f4903abfdc7b74488",
      x"8b4cf18e273ddc06fd6ab2a09dbafc20830a90ac1401a168aec5e24375b8415e",
      x"775c98c545bc10a7643efbd4f59bd3ffe193623582cf5c72c4f4be7c5f286429",
      x"eb2bf3d488d7b2230917076cf17b08bac61781def67ac31915dda6939ad1ca55",
      x"13b21e1882b0ee0ea4519fe1c0175ed425ed872c50e0eebe7c88c3072d51aff9",
      x"06e28fad1e3e25b57e2b337bc05420330d86e958bc405ce708b14e55e81a60e5",
      x"185d64362c39f3888f9250121f922974e3f06957eb5ae50a94fcf20054e2b780",
      x"52347f18bc5e5c0bc95dfabe08bfd5ad33b6a6596fc7ef44edf1231e8ca45d9d",
      x"c3c98483b2d6b5295f070751ed776fe72422234fed5014622b6d65a2f74e8fdb",
      x"4a9fdb977e8f334a567b2a2fcf0a4c6ca519f5c296162787332eeac98b05bdde",
      x"523c1a36f6d9da00ff7ed50771b237a97eb3e1b21bba99231aef92747e2783bb",
      x"eab0a2e44c2ad627ed536e19c8642e0e2a1aedb21f0799a03c0237edc3c06fb8",
      x"c4e3dce074d330295f4e979d164f2ecfce639fe357c4ae6ccf544d6d23eeee4d",
      x"5b966910ab802553e995d27de677d7e6d7ada7ee77ace0eb051566e16df73153",
      x"f72f3caeaa0096f19771c2353dd8f7eb0b6a09b2ccc99a7a7abe1319196d6747",
      x"164ce16380f657f7d4841219f897b98e71c5da569033cb1c1580d9019148c2ab",
      x"7b31cabc4b5fab9bdafc8fe17ca9080c7285eb6198959b9406d75f0488fe96be",
      x"e7c7ed870973819b8cc87cd102c9339a7e726918acd599c660a924f1cf52b08b",
      x"51958c2777ff2dfbc3e776588f56920c37b9331807a51f56097316e856f5ac27",
      x"617d6d6437680f44e5cf6d34505361d7511d685f9a43fac5da6816423e22e927",
      x"b9a7219143b011243d1c2d4bbde7fe5842094c1a17a14c8d960210f88992769b",
      x"671210a1ce176f7ccbd24ac449c029bad5fd4ea2f7299baead6f15ec1cd0cc1a",
      x"53c5f2d7154a4ff2b91088aebe5d7c00933fda5cd33fff49b8ab2ea0205d3d3c",
      x"cb729b32681cbb1adaa356f7bfcf381ec1db95d3787d2b2afad3ce0fd6744e23",
      x"a61c36c30d8f0974034d4a5c15183a3337ef91c3eb1239c180826389dcb75648",
      x"530bc2d3cbbe3d2a8a6143ce4f79983faf0c735ce8515b01bf609858e01205f7",
      x"07e27f5322e0d35ba6c743b0a238d59700c62f507c84b799dc780e0e29f7ae1e",
      x"4689f6fd287619443ee2abcecadfaf451d526b2d77606ef5b85b6869cb183f8a",
      x"12138ae01baf0e47d56b57a39af7841fb73f9c98f7c41e88d6eaa68699e3513f",
      x"84dc707d7b1a04346868bca5a1cb3b8feeafa0f9461e1ae8ae3dc40f1b7ad07f",
      x"aa242d21f5e6ad660de684ac33af130742919312296bac3878eedd2e2a1bd81e",
      x"ebbd978f5bd8ecbd57c767001c2bcda7a1e1085ff9141727338a55e9b14dd98f",
      x"5a2c10765d2a1cff7e0faf1c8e33139fdd0656a504fc6b4db188afa88875bc1f",
      x"810d23196b08fa9467efa11fc471aa7a1cc2851cf8410ba592d90dc47d2565a9",
      x"9c13a85d30eaa252ded4f16f95fa693b672c41ea9c6bf5b2d2b12a193b0e52c9",
      x"c604d95938a5969ca6e3132917ca5e404a853ad412f45b2c6478f6d57050da34",
      x"ca12cf14c12cc8d30257eacdbcb82ce325fbbea63da92e3dccd402ef7ebea6cb",
      x"80c0a3ee391446eaf15354bb56d1392b9b4a2c89e5fe460ec767949238081957",
      x"283aa63f5a7e64934ff0559c4fd260871001a1f4468a6d7cb93e5f5dca2efa99",
      x"3d152004a376d1252cff41e2e801f3c537203d0d4a07b7eb3392841a58c3c4b9",
      x"f71bf7efbcb96e1a0fdd4876c2a2d17e97af7f2fbc8044798b7c01f467b4cac0",
      x"82ae2b412b1e1736bf2b7663dc2774af61f375aa099ef115ab252c77ab623c8b",
      x"b291eed4d2ac42749918cf1c09aecaf589fb1ea10c45b2e7c336ebd4efd30ed4",
      x"5399cd0b0e12112cf8e841c7a176d60e3ad1552600068004bc074fb3ee0c3cd4",
      x"ddf090e4d8549bf33cd00d813a612bfb0d89f1fa6718af9e73a0a5affff50b3f",
      x"02ef3fe16a5f610f92619328ff65b05c9d8cca73be00dbccff737ff6f1405939",
      x"17a7490cff7a827a4324f2750fa9975d57bfb8b00a678eb8c06101ad1ea3e967",
      x"597047bf05a046d26e2d6362db77f82d2eb6f2ec14e34765a0e480531ea0742e",
      x"d6318652d074f38259fe26b19ad669fa91ee9cc93eeabc907955bb2724f412bd",
      x"923aa4f21cef7fb30372990b363731b884d358a3259418e94823837640618278",
      x"2f84484d286062bd89efb80abc1c402921e6dbcac7ac5ce1e8a171d692421c1f",
      x"b603f746ab35daa5b0129105e72297d50c5b6d12efc7e4a3da461b4994cafe47",
      x"dcbd650946e224fd82f62378da46f870a62e4c34c46156e3ec73c67d63253206",
      x"9ac7930813d656049b6863789db1f2c97f6e9411a6114e0107ed68c41ba9f575",
      x"b40f78db6661f930c72f1e9f1fa84fd859b564c32ce3c64a337c3f16de106734",
      x"db719e5edfe8651ca10e34e090f1f36140e34a283e2b75a22c55b87025cfc57d",
      x"0a23cc3045b72e1350581ebeecde5c3d31c4fbb726becaec9c0131defcddc59f",
      x"0164d39dc54735bbc6a576bb9b3ef3705549d59282e5469487695c864dfe17a4",
      x"e43b3d6e3b1ad7a3c5b3e5b4ef0b2f260df01d2ea4dd183010fddf535695dd75",
      x"31eed53429b0c7ee2a6facf4cd995f120840c261d70acc7d9999294943f4e99c",
      x"45876b7e6a82bd4873e8e81025edc3d333a15684303d70a7b58ae446b35a1608",
      x"3f5afd9245c29629beab9c56a1e8830231135a42d9083596f78ab5078bd5bf63",
      x"bdb9b4f94faddde0de9ee0b0a6261a074f62a4bc66cf79c4abf03ab3514c97bc",
      x"4c465e688d38d4e855396c8661ed368915e001a1c1a6b512a3854c878ca18d41",
      x"886481ca540d769a519e8d5cc0333087feda78e4b2e23909e07ac3f024930325",
      x"5472575edaf265a33fb6aa3bdaacf4c52fb95722ed02da2ddb3d26c2bdf12be7"
    ),
    (
      x"65a042f2a90f45f47dab8b7c5ec80dc55c0ac290abc9430354687513f221971f",
      x"09eea9be5b01ab75c47677eb2026bf06000d9ac7de3b87a78632be671d103dfc",
      x"6b3637f58626212ecddbb306318f6e856ca2e282b0614b159c799c8f52540a2e",
      x"95b828e9bb9ec1d85985e13d2b7504debe050f96149518ec775b2cd193d26a64",
      x"7e5b0781de90a56df9695ecf4ae5b2841e4d43a568e8a259f3b0de85dd0c4eb3",
      x"5083017950344837d844c04750045a97379f107ac27815d1f48794d5456517b1",
      x"dd2a1de3ca0a657b3760f0c9f705cb8db1590342ec6b6c9731b5df21f334317f",
      x"8db6eeae5ad573d84501d45040d94a827d215956037ed9b3fa3cd06a05a5fc63",
      x"1c8b42c26d5d928c86ea40d5b55d8307038dae2628e14f9f7ca2a8720d9df784",
      x"cfdcbae3103c0a19e571f3ce13f0ce04728225bcbd7aaa6541db0bfd28253d76",
      x"ec67c02569dafb688ef59030f5c7c92f47314756ff9bd853671a96098b848ea3",
      x"cefae6df3152ebbda506e875c84cb4463fee032c913e7f9d875ea0fa4b65bd89",
      x"498c7a90e0809899be81533ba8e625ad0e40e645d2b11ab4cc4afd1f7a61a678",
      x"8b360f59b96c76d1697d23970f7140ab562c54c4c0530fe964b3891c8f1010bf",
      x"644e8d6c8e313daf4f7c4b8172f205412bde3c1d18249271574a0d30fa5e2075",
      x"73f15803c5dc057f0cbad45124c64bef7c35ea6e36b07baf867a5d9ed48aeba7",
      x"2610c8da6c78eb55dd806399d0894c99e951740b67562d0812c9e881f0403613",
      x"db404d8282a75b0ce38d96dcecbfa3b98e792f048df5b59f329ece2155656d0b",
      x"ca0fc91c19093050c6f482882273ac75694ee8ef6496e04310821335a494ad2a",
      x"de9aa68aa2b4a6daa388f479750b2c24bd52f41233da42be4f8c69a5aae1f2a2",
      x"965e7e1fa8faabfd965b1c993225866db04bb00cb3b0d2aac4ab078bb9e20d7f",
      x"90c928e67c8628e15637e0f57763a166fe59331e1c54f8083cd28b5127c09af1",
      x"85c4951229b9eecf49971b0ea675cc50b1531d8de8825b0c3f33a1171f5ecaa9",
      x"32bcfa27372dba9420cbc30fa3b5f607c7496c2f72e916e9d8cd2154a62bcbe8",
      x"94808899cfb1d7513e9a83b104c316b7a0100ec2f72c6b923fa70f8d24c13d87",
      x"b3c29bd02652622831034933b844b1a79e2312299a340246a731682d9923ac46",
      x"8be8c70dd5315348f6ce24da4a6e1bc3ac7062979502ae5550cc733dcbdf1b1e",
      x"095fdf637c0fc3660e4b20dcc0627c28d0ea755b2fabc872cf07b3a94050276d",
      x"4d9050e549d5f47eaccf9d057c328e7f30b7b6a921e4517917578782b3b16003",
      x"b5a14ee3dedf43084e7449d4ab42ef5fc0e8e285775bf7126b211381003e4f4e",
      x"a38cddf68ad27c17899fe8bddcf5b5415390cf2a7cafc8187c38e60e5df4864b",
      x"1b803e5a9a745e62a01aef47bbfc43543b76946c7f5b1f2d6d54818999340494",
      x"0544c009e8f63881f3ea58b82478e028959e590e292684fc8e23203075369552",
      x"b17282a6747062d81fa3447796234261dc7cf4ef3f626852f8e34abc4bc56168",
      x"b8067987d49546bbe0ad2ee4992566f1fc1f48514eb3a24fbf2193e7c2fae942",
      x"fb014a7e9c6e9cdb5eb1a00f41f859f5dc763acd1995604f5f12a6dc76d68e24",
      x"dacb8f3fd8e03a6d0f4a5952312925ce9c7a39c52dc298611fdf80af57262df3",
      x"76b17b2d5561c139dbcb6a9705ebe78a2bec20fd041be70fda4f130360e743c5",
      x"3bc4f17f07bdc990f542ccd635e2aa5fa9c9bed0ceceaf553a2780787a331ee0",
      x"d23f689153d711500f671af5c210a1b9e38e7de67b5d0092cb2b9a1a0e953c80",
      x"e5a651c64352fa62daaa27aa975b804fbb32366d51c78546fa7e2ba9cd2f153a",
      x"eb77c3fb97f5ee09660841bb238543ced954320f04d58b0adb5e8afb63cacc46",
      x"f5a7edab7ae3408ce482e614a9be18a248b69c658244485e9b69f0f7fda35957",
      x"0c2b9cc2e215cff30614c014cfa8dfd876b9be737fd5bdf8206572cc3af7efe6",
      x"e813d8ca66a9caf7d06673d7633e337855df2b210659fb2923176d892e9b8183",
      x"b3398da112d28d7980b125bf041b9b5a071e2f69a94895e5aee011a7e2c5adb6",
      x"6cc9c3d00bec038d493adb58048bfc7096fe8cf958a63a4cdb75da07ad75a9f7",
      x"a309abfe11ed7c3db5c553cfdb27c713d3011490f3e2cd37a6647ac44b43cbfc",
      x"14bc588ff8b735aac8fb8343a4a8ebe5cbff2ba706829e6b9efa34bff311eb0d",
      x"7cb84ed7e233547d8d239a738acfaa364360d1fe1cddd6f335c116ad4629e31e",
      x"b24df54de47dcd3ef40318b99ced01ad9307c73fec517510b363fc06b1f15044",
      x"9f5b7de4b3aaca2699d4b7056c29d42cc0d24ff6b8f87e89a73a8254a3524b4b",
      x"050492e6d2c6f1bac9591485c95ecafe578104dbf53c484db0605a3ca0ed845d",
      x"516d5132e9b08539939c50f5bdc30d4850d503b4e3389a93c3ca1c9c333f8edd",
      x"766d62a22b354b20dab52d00ac65106aff59c814905aedc4da32b59298d65a4f",
      x"f8ac0080d2f3fba50d635c11946dff48b9c75a7ce6b874695e4934c04ad7d082",
      x"cfbb9225c5f2e04d095de8475d127666ed5085dc325e6a53eabc23707cf2449a",
      x"85b8db23d367f0b9c944f9928ec40ccd1d2e495616b18107652f1b6955ec70e6",
      x"e229f68370e70a3006a17500026816c2374c3d2b2e23d249e5e76c0741049914",
      x"2d26334d03a61a01d25956b9adcee6c4c0e8acbe95af42db5bd8488f868e217b",
      x"760d91f163e69e868905e94de06af87614bd49f7444a64d6c98a3e002c169331",
      x"2e903f11ce4e2a808f4698d0b824993dc0a061c70d6a1e6dd62ad1330b3484eb",
      x"bf412f9b22199e575a2fac99da07b9d2f0fa6bfe68d92fd9d9a6d471a4eae566",
      x"948842895621de12adc320921655e81847b55a64196f8bda059f74e7f51e466c",
      x"bde462b3161b32b265003cf21a21e23d60198d9a5d3867964efe208a0992b3a0",
      x"d6c028e4e4f8a72fbd5ce5b3c43be5e7f856fbfcac5648ee398ee6ded5695799",
      x"4451e53785a45b6d2a32d02789ebcc96bf4083dfd6091c257b90e3cdc14b4fd7",
      x"1459111682a53c31c089acdbf0d6fb175c2ca42f68815ff0ecdf9b83f51cc563",
      x"1ac5556b47445a3122316af5fa1edd9500a18c66640a0d622d08b9b26e592df9",
      x"5e14e334553469906c61229569835e5bba55bded09ced77a1217872b4c1d8982",
      x"0e367e3317383d29cf011ef0ffe54869b817c8a810fedf31e06a66383b8c5465",
      x"41eb654932cd741c1c1135e4e021cdebfc8452e2a9b478eed6c3c035a1532fe1",
      x"a1b8060c14fd9c4dba272204ce8add0d29a754e78dacf64e0c8a81fc18a808ce",
      x"242e76202182c359696b5ad817482d74a9511af6960588d2a3bb1fcb416a3f50",
      x"72b8532ed16bd8faba654a1c4f5c47b9f0fe63c9ac35215b42e04cea21773b7b",
      x"52810f1a35c9ef7506e746680301428fb4524afff879759ce6057ac796ab7282",
      x"824ed3c0cbcba87945d5941cc3fdb6042fd62373fcb8fa83f81903cef73ff9cd",
      x"a118ea99d9d44e880ff1e8bcaece6e427ea90f2ab9914ca8d38aa06371281902",
      x"98b4c392fc8428146c2115b223a8035f54022ddfade03ed20508529694823ca1",
      x"e532124335f39b41c5b9d0f12a409312bc72502f11f1890be6e4f83f68c3f96d",
      x"05f1d2827b76688454187e9fda73f098bc7488d2256b58be5986960ac4505f47",
      x"033a0581e6e7ceee24d11baf5117ace7de7b5732bba3d1685d3a9f45ca71ddf8",
      x"3357c47ed63fe8be78390ba98e5be15134e3fe006519c2f7c3ff29c90a0864a7",
      x"a4c612b99c1d69360c569970ce15d802693d96134de55067b8e18719e05b76cc",
      x"7b220faa093a72dd6057b0146c43b837aee6f3c716761a8b1d1e2e273fe6f6c1",
      x"0727887a30d0379e9ce13a73ea68eb2e965f6676857ec5dbe9e772ece721e213",
      x"aef7133cad950410e9a68b6bc28f92e4f3f2ca274b16a5551a78ce10b40c702d",
      x"63140d60e1bc01f06c0fef193618a22f90fed0f71bc700d60e908fe2701ea9a7",
      x"f83db716498653ddae20e3bf9af612e2c219258749fbc014d04f1354f898542e",
      x"765ee305dfbfe212c457a054d363ee8ab36bdc54650fb0a2382b3f693087bc39",
      x"621068eb57e0cf5881b072b803d1acdabb1458558a131b03600e8e85bd0c6e34",
      x"a96789582737c879d11454eb1eb231a831364216de0e4906f20cf69bcd14a578",
      x"0f8647f4eac6bc3c926a9a4526ad9523b71d70c5d67c66ed43dba274b3db4861",
      x"2c88ede95a88f015f8b9a3335b5e8af07d9cf6c5e7ed9f407bb61dafc47c4afa",
      x"20e8d6f6556ce5031cbba7c7d6d2e8d4f7e738fbb69b00ead9ec33da4582bbb1",
      x"5fcc15ab2f71a5f00ab36b7795d15aca4cd9ba0900f1ef606407fa3969faa454",
      x"7f5db6b7b746a06d6c1c504400cc0127955ba318246c27484148a11baa58bba1",
      x"3aa013a82c3ffa55c694aed0cd5419e2d4a98a5d22dd4c17a402eb8ac1c1873c",
      x"a3dd4eb021d76337454fc5ec45800ee6a89a46fa9a5711fe6cc11435484def0a",
      x"52848412505648bad24f779436465a1967ce19b1e882cfafd5b355a646112541",
      x"eaeb124797f7904ec5c2d2e2d5e29fcdb0cdcd61ad5bb44b676af92e693c42cf",
      x"6d0d2b9c98fa5660ed594804e607cb6d60ab3f228d61b52cdbfe4f10c6cb2492",
      x"d4aff7738a4d004f988efacbb936bcb3f5258c03c216c3db14909664263fa403",
      x"cd91018be6dad2161a67c7fac5a2ce47cf3c714b98e98ea7de64a1f60fc991a1",
      x"fed51aecf9330e7ae0dfff25c20b1bede15b41a3e7ee3f96f536140ce566497d",
      x"b5b3804a3fc7ccedf869d30aabe8045e8020b60988e7f77b532ab3fbc8e8a1bc",
      x"1477736e53018a5c3152119d9f006539f093dc7cb63a89006a2247bee321f3b7",
      x"509bae85b91dc401cc1047b75fba26f635454937bf9b08139e9d014d95e5bd15",
      x"9d171ad035ec2dae14b7d7e1c234100ae9474642e6b6d574dcecc14abba19f67",
      x"cb6894828e59f5f2a5a8151af6c5ddde4e559690e47c539d31c76b6a96da56b1",
      x"78bb51c7ace2c94e337ad7ece4ddd5bf031562513f9cd4e6fbae5bc14d4bb05d",
      x"d930a46c1d0e4cebc8074845e4276098ce05ea95e27403d00fb948dbce332d7d",
      x"dbebed22961bdfdf9ad753934c5bb6b54a5fd17edb5b18ee500d8fff84da7264",
      x"398ff83f79e0d4a5410abcfd42025611389fe11fd6fdcd7eb9af71f390e0cd09",
      x"9a96dd4588a0bd0ae21288e06d29694994f4cb4a8dc8956f382b0a55310df32d",
      x"e337555988c7eef60318b725b03cad90c597a7279e5d0c7077c53d5ffdb36916",
      x"a0fdf10eb6ed315a94ce8759555e84b1633d6f00688842da120df6a894751d6b",
      x"bf70c5544073e6d1473ec086e8772d06b516ce4294981f44d14c828ee33aba39",
      x"562451d6704039b7939f1e4d8572392a921be8c0a625aee7f86c8ea996a97e93",
      x"2dc08d9c38199ab558522e63eca5cc247a3246da0e1ea567620c5ef5686bf0d3",
      x"783d0372da69a09084e18fe1c4f8a1618960122bbc3af8bf508c3048a834e50f",
      x"982180ad4a97a32914e03244f89f88434d80c467c2b0109e25da07f6eb5010f8",
      x"2f16767e16395ee93618829df595e2ef65f39d4918d235e596a3217246f3fc97",
      x"b9d0756ebac9b08e9ce0a43db891e9eea1b459196ca109139f4d2defc622f833",
      x"8bfa19d8c14d5d2f3dbe4510e2d6ff6d8b2f76c59ca39fff3f1ec87676325001",
      x"20af2f4e912b3bc8d5e3999aa439ac5e2a7081a904f2548ca36e1c1b5a0d74f8",
      x"ccba1bf96dd8779120a49f1a16c03ffd24dd0fbafb1b6838a778f4551ecbcc53",
      x"262889830487fd183beae10c025130d52b111371d620ffb9b230cf6b16bec129",
      x"ee9da97bac0778802bef5631bfe4e3c3844c35e9702989a5651aca18e89b6dc1",
      x"02a16184a3fde321898d01e21c08e253c3de00d6ac3c92a73a657e9539c726db",
      x"a7ba948a5ed489c708315874144604c17a96c7bce816c6d13554a28ea2ea41e3",
      x"239bbb3ee3abc572091a5da3dc5f1614a41bffd8b541b3574d30e1e2e520802b",
      x"9476030cf38d28162c907b6cb800f1fbc93a641dd0cbd3bf9d64537380c72cb8",
      x"cf0a81f045740493cc905d346dfd531ba0ca7c2a5c3029b5ca4995d7bc4b55f7",
      x"c7b88842ead756dde6ab8fedcb7d6a6d3cb451c161662e3b31bed61f0bee1c69",
      x"913c7eefc7a144762bf21c0027927b1e7612f906cbf3d40644b0542516b31499",
      x"8bc8f514129db81b7bccddbb19ee6fedc45bdc83ee373ceec99f44e8fff536d4",
      x"6b54732781af3e01baff3f28d6fbe79ba52a7eae22ec338d920630a058a8c1b5",
      x"12142cd08d531a1b3c7468a3f266d72f294614467745dfffdbc7d531f2fdff07",
      x"9bf0eaaffefe822402604eb5f78b2a3d78559121d35ffd59d0fec600aa4d683e",
      x"2ac9beb28c2268259715ac2b999df762aafd5edc16450fc2644e4c7a976354d2",
      x"4c49beedca6659ab3ac5180143bf876822a63d5dd07b12c66aafe63301ede668",
      x"3800d023f380bbc8b29d5f819261942d5023215081fda37cf5baeb6f1e2b2a10",
      x"a47d4c10e354af5f9bf65ec33bb9f5ed182061356b717de589d96099391283fb",
      x"ceaa2c8b6db4f434fadd4032d34440f88936443f6d3a53dc1975c72ad87e6def",
      x"b0334c80d2b3f2c9c90f58fbac8cc155b6c3573aa1522fd79cfff29222e6ea87",
      x"05fa62f3c1b9d3a5ab04a58e766478e2ee7ec83c6395935de46152b699dcf7f2",
      x"56dd61bf2737f8d44b57742442ae0e709dd2461b754d01dd7eb90fe40d372c3f",
      x"6cd8803e482c0698e8a9eefe21327061dbc020c415b8b89d511c921d87a2c7e6",
      x"19224445a7605f392cd301968543b248ddea8bdd18c938f3367b2a4678738bde",
      x"1fb7be7d0555fd82709bb631628424397b104d891e1d4e3d26cd74423c01ea9c",
      x"3b35ae1f1d6326873e06ff0e191678692d434680f9aac476196bd7b05446cecd",
      x"41a999a251adbb19cc9aef43c8933f770c6a6085a6c44879a682247d5fc88962",
      x"38b5e495d37d333ba17d21614510a462c53e82fe0cf7bbf9afd9e100d694c55a",
      x"547a7d904efbbe8861b8e86e93d2ae1345daa433fa1997b55aad69fef965576b",
      x"e3b3a21f2382ee4a8dbc2788bc805e3dc2d1151590fd27096a38aa60210883d3",
      x"7a2205f3d11e36de9b11a739bc380f0752ce1580c4a94c5439ece86e844d2f31",
      x"c368d31e601afd753bb3aff2eacf14ff93732639810d22154d137f2d80346eba",
      x"47c3d47bd663c5a1283979d5d22f9c5cd949104f12ef45a789e95b9a171def0a",
      x"fe36daa8d89f5d5aa2c1ab5b46d181b7f5da5955970b1d9f730d127214bcb56c",
      x"8b20f9a11fb9cad6c22a0f6da8f75bd66da22fcf7661ff0fe6093086612936e3",
      x"6f10ef452f7765b8eeacbdbc574a9064064e95613eb88209aa201da72eeea600",
      x"ccf1ee2077a81c2ad63b0e67598f19eb586c098074b8c8575efb005578a5aed7",
      x"1e6f40db37b3987af66926e1722a87f2233c7b21efd9461ee6bb069e24040547",
      x"2e4ee38a732026434c527c64ddea35250e38866a06c640b22e833dd7b57fe016",
      x"c1316a12f260fbb6f40cb8a83645590d1610e6d03969a6b5b05049f03a65caa5",
      x"64581ba4a6c6471fca94cd93e16953a9ff4993aab1547581c2a57ec51e53d2f0",
      x"54b1772fee140092d3e43a2d50114c0a7548ae4d051f479ece14cddb0630e587",
      x"df6e3185a386bb0fdb5becba9437baac9c43f5943b01a74e49a4b4af0ba81f7e",
      x"07453a01a680a7bd7c0045cc9fc78d11b6058fe7fc4fb3b02e5340123c4de996",
      x"82359184b96fecfb7c7cd43fd629a14a6c021ffca1138d471e779526eb6d1e1e",
      x"17acc653edb3ebaa9ff171005936f9b6da17947b4f2b59daf00decbf7fc9b74a",
      x"2c7986238628b38659e92a185a1559115f15166d271ce3401a161ba4491890cb",
      x"8c7d3b9372e72fe1862680aac3e64c2c88c3008f8e8615cd9858e2e2105c40ac",
      x"1e92406bbf604bad20ec44b4d0ff2a1de1aaa5d8c5ad4594275a0c6f9cbe2f08",
      x"903d367a7f06bdf605e0dfacc0c615f5be03e1988b6e15ec6225e3cf390294f9",
      x"2f552d1518f21732d17aeba053b1f6c7b272240df04c62db40dc002860aeb78a",
      x"531e77094c44c11c6bf79033e93e090b5af9ffc8992e9a777d5697b37efc259e",
      x"418f41db83c25b9a066edb588cf96196655ea608868e6cb8fda268d4d048e952",
      x"81a796ab0b5795133fe67a6d39781baf8dd51957328013285d774e499c92a8be",
      x"1d87b9caf40b625defc6c0b518045cae9ee4d952562082f4470dce5c497b4b08",
      x"6ff272555cc417c08f312aca907c8354337a6c6ae00794458ce68042aae2da55",
      x"f6313171fd32bd26c16a6095a3059d599c582c41de3c24d4998a51a6b19ab014",
      x"4cc8a95ee9f95b87615e823899b8f8b787a0f3c579e64bfc857db44896c41a86",
      x"c2ce7668ad6d9e3c6620aacedafe4acf9f49e78fccd1aff12037b842ea33bcae",
      x"f33b06074d7a92b162cc20db11d205673e64d3af484186c64a561006cb864cdd",
      x"564684c34501ad4e8a6c9a591850acec9a61d4c8dae8d5b0a6fb5e16c9911b21",
      x"da3856ce5beb71898556d66a8566d09af72093284d14717ce3177d9220a4f8d5",
      x"ae1f06d27de821c8ad7d05f3dcc607e7ef7c21419a036e614dd68bc8423cd4e1",
      x"c2e672d70c7b2cde637bc8e3ec8940441eb2623bb2a5bc9c64f87acc745163f3",
      x"b089f69c2b5e59b901fc8c42c34253a61a5cbc9b5615f5ff138eff5f74829387",
      x"14f9d99e152d99aa5c26fe4ffd3d4f9490c23f044109179023ab115b541d27e9",
      x"db769886aec47b2e8db50b92e18f4cf56c0e2d69d689c204281680be628d5d8c",
      x"c4ac150197c572e8aa40336927428edae8935fa103da21a90315f4de9f80a375",
      x"f5ec236d11604dffae1b5e3cc11cf11d7c97bc578d3e7aa378c26aa07a055dac",
      x"594d541ecb83db3a35df36ab1d7a1ca82cdf005c724bc9b1610b6d603f619630",
      x"a4a78bd281f88a6dc2ba39b5b83132037a7cca1f0efff67ac8954524aa6d3101",
      x"5c5e1322fdd9e360f226b38b0a99cf53c83ded73b2cae2291a7b0d7d594c83b3",
      x"7890cd68a0c64991d3ad5d776e703ee4901a355dc18f9e20aae54883dbbc9dd1",
      x"927c07b0171c94e3a5811b17185b60ffde23a3b6a2292e3b9d40d67b19fef25b",
      x"f8e32ac448409a758ca53560f0aea7f92ac416c89474b8e1f20fdf58ad62e880",
      x"8fdb8dfc06c87d049d6dafcf5b9202e4251f310e68d8162c337aa38294565142",
      x"cbfca4350625e8fa2c4c19f1409dc31faa46312f06d9990ff37fc7b0c6d0637d",
      x"cf00abcd2c658f8d43030790e2b7cd87b23e6de437d974ebbf52d66c250a52d9",
      x"6284a063c262ef861f6e34a55a962e9a3ce5219617f59ad21e9b9897a8d26bbf",
      x"af0647a449c6aa2fd4a59ea7dc9bc3832aa0368dba48b6b60f2eeca817775ea3",
      x"6ef0012fea78a2336d6fc56a6c867a74584bda4acdc0caade83393faccec7b1b",
      x"be400280fce6a343ab871aebdd962336e7c5bb5fde853d593f3727812dec7330",
      x"cf09b981970a50f1874556eb6dcb0a31b3e400c8d69e9de894f9274187cc9a8e",
      x"2163f76a93c022ef935c28e04b48f5fa7b924dfd641c7a79fa2d6149a929012f",
      x"5758e7ce0e856146c69b4bc03f0039e6b57ba206958bb2bb0eb09c3f40781004",
      x"5c817e8bf4d4d677e5a9cfe6c0bad254ccac5f3952246aa1a473119945f37cd3",
      x"eb9aba2e9fc426227cca13bd89664d369d47f8bc0677fb1f4d86adbe02122ac3",
      x"465923cba1719a70b77f82122301bd81a0f4db975dd687605ce8eda72b957eb6",
      x"30826d8a1410f1c6ba5b30a338a0b68a3735f20e2520f62bc5f8dabd68767ab9",
      x"d5324ed48a30beac1326057e65db047a93af6a53f9900b2e0a68369e6ce27724",
      x"99652a14f31cbba33fd7109fceaca081919be1d35047c6a25c6276fd6b27ad83",
      x"da8eab12f2ce1bf4fca5e80989ff39214e97db861120341eccd44b949f2b6057",
      x"88ebce5cdba2959717df644344479cb2f6d6c6b3cae2a01bc70e10a25b6ef60e",
      x"6803cc570ae3947ef85efceda0597b0a0e4d6b46c14261ec0bc035c3cdc66539",
      x"f62650f00a81db1840dddbe776ef124fe5f36b0c09a1553e17688dfe4485dec5",
      x"947bf00132e7b6ede5a6d349bf5cab016f633bda7f9a6ab6768f8065e3961fc5",
      x"1c77dec7a6ac4d35e31a3e6dac3a9d1a0558ece1f7d569f52f90abbb606a0cf4",
      x"08d3ce35cc95843a6c7629474ccfc18677bea5a676458cc0ff4ea9304ac8216b",
      x"1c68774e8779d3747c5c942ff0778fe415dccca5ce88459da216257f849691cd",
      x"6c84e0ea99b6bc7c6f11273ee0486827947470b8011af062704418ea9cce06b7",
      x"9994bc8dad9fb97f19651fdd3f5de070535cd8a6d75d33a22b9a35826eaaa570",
      x"d1d19903446dd113e875ca025a16286e60f8dc2fff4ac19911d66977cb33b979",
      x"cdc76825e1c87a74a4c722a72209042534c17b1c0d2cb182df2c5555798038ae",
      x"96d91249d856623aaf504fc509fea74664234ffbcbc8eb4d568e9857760b0a02",
      x"faee1db3ffc2d2686dbe9b6db2a1d41fd62f079dab30039514813bdcc0e3974a",
      x"2240ab2285ce0b8121a7067efeb4eb44f9ab5c9f8cc68c97b13a2fafe61c0378",
      x"96a7766c2935fa8ed2609c4177ff035dc4c349530d4ae93234d32c445c9d648b",
      x"9da3c935858032d67e0a8353a097c7993cc4986226805b60834ec220ebd9529b",
      x"7e9ec54d1a8991f384c2968eaa33111cb6a9ae83213e5f3ff7ed1a539d2e6b74",
      x"fb37b035b24a1fd0752a345a83e3794fa4e5215f7aedb1b4c81babe2b78b17d0",
      x"c9356efbdc2b3af4e8c364ceb19323d59ce93a6ec555271e017b4d21e9eef2a2",
      x"53665e4bda1ceaf85905a8739ca7191e5f28cec958eeaa736a431bd217ba9fe3",
      x"a81d260a229da47f2cf0e6b898f5c0e6231a2b6cba289b0f66ff89f48480c90a",
      x"b717fdc6ceecb5aa0404c476757363646cb18b0d9f87d51b16a457998f9d28f0",
      x"8ebdf893f98fe6d726883e782b8d758214a1cc0237a6df6e42d2cf18b7193e83",
      x"517829221d2a64c639a1cc4c025652f320da35761cb9b208857b21f7025fa571",
      x"acab5828f3436316c555e9955482ca402828a0e54a3a1dea3259ec2136d1e3d1",
      x"a44c05b31e6d60cb56f773dc228c52c9966717c9e7c9a671e6f8b071f144f69a",
      x"d6e14c7b23c3b69f2d6ff49c09e76659378215bf9912d62cd2dbe4e48c3384c4",
      x"0523c3a258c5461e88daac7d0b4604d8f05c1a08b8abe63cac51a050f444e36f",
      x"42335e9b092287e211edc85d287d5beb53c438505f4f64488f0d54dfd568373f",
      x"6f6566d330b70bd8d6684a5b6ec241cd1190d1a38d8f12ab41d4beb939b6a375",
      x"4ea36618403a7156cc6943b67b7f20b33f4410ee6b44272f59a0f6bdd0d00daf",
      x"061605c9178258d7c770d6484a06f62a1affdd2b146149a61df6bbabf87751b9",
      x"b02f2e72169e148050099dcda484200dac12ca7992a2f93426b836d8fc4d1185",
      x"6e4cc026e08f3a5d1a1d1724aa5b285812835a6d10add001efef7cae7b525963",
      x"69ed0b1df238845b14ada1fbb3b78250c3a7626f798308b1379ee2f8c0f97b33",
      x"8d68b8ecc545f8303ceef27db171122053e8fa79dd2535b17cf931ecefbd9387",
      x"1654fdd17388114018fc6deeb680dfa6c1d1bab982e91e1d5f690647222bd829",
      x"db9bbb343362a73c8b58815f3183275422b1b5cbe11fc8ad6ccc329f12cebead"
    ),
    (
      x"ca88a3f31f90876e24522ad0d1f4489bef167ddcf9ce2c23bdef3cf0af2127f7",
      x"cf678edefa888cf8918a7459c69e89f10a77bef45325fff4977b01afdc40e884",
      x"60754132e1aa4dba3007f5932c4fcade84cd28c15289970fb441f7334eeb0933",
      x"fb854b7f7ef4d32561cf0804f1a31a4a3acac8524fe56c0df8f1c46ac70d06f4",
      x"26a6fc35e167d9bdec2d3afe97ef1f532a636024f1f69a380238e7dffdb2f763",
      x"d57ee32d065ce346ee1ab71debeb522d8c001ddcdb6a90fa240cb294159778dc",
      x"84ac7811b5a508e4b3aee3598c537267a01cb34b05a26910b5c4b36ee406ded2",
      x"8a0759213692958790d536c709a60fe292b9e09c7c0e103af27808b03df43b70",
      x"0b39586bd81fdf29ace1f206522282b2206d9e61b5836c4d22669f318ae0e767",
      x"3e0bee509f49c8b80a625705366192c888a0ab1932477f8fccdfb0aef2fc79cd",
      x"6f9eab3c6ab0d98f0e52fae35312919fa362711d63d21985a1a84cce00fa115f",
      x"93ca254ec36c113bdf2daa10663d61f923979531e85560bc7c7202abbc1698f9",
      x"d160b08a9df83a2bfc5460d215670f500f126d92b02d1ceb5d719f482cb84ed6",
      x"57cfe300b680f8b2070469c52bc65749e042ed60d305e12c54df1dc0398ff65f",
      x"f932bee76b4d03d46d16fe78eec25cc84809ec7803fae0e5e4272d7131e50cef",
      x"5af23072c9f764ce70cfa6a8e7b7924912642a21e5c1ad6b90db26be94347a69",
      x"6204a39d7c661a338dd4fa34084c3130fd4b3ed820c7ea93e785e39904039919",
      x"2178c2cd6caa473805feefa50c4963f62f5a2f4be0db9aa444e666e2e49654f8",
      x"a3efe96d13381cca8416245035bf5f79f3d2897b559ecfd5f4982f7ceeeb7c93",
      x"1b4efcf8ce4befa287e63e74c1480683e05a37f176f21c2af08afc73bd07bfcf",
      x"119b1defbeed38554c0cc653d68651cf26bc39dcdf68fdf36e5a944c68dfb012",
      x"dd16b36bec006823c96b2201c34c31bd22c4875e9d7b34eaaab9f6d2f59a69d8",
      x"fb0eaad606135b3ce1325bc34d0098423eaf8feaf160479b460a30369de206bd",
      x"c79011c6334e1dc0830887c98fe62ec8183ca99112b79e3ce348d666dfc79bee",
      x"f1f0e81680efd3982456ebd0045326d8c45b2a37b7325f528cdc9abf187e5a8f",
      x"76834e959fc41d453b484f6ce4ac7f35d68f9b548c970b6a5635c7ff26528a39",
      x"4dd18eee8048a030ca3e24dbf6569a180eb96288bfdad20916eb20e486370b51",
      x"8830e7fa8a968606805508e933e77eeb1a2680e5aafe4e5cb4499d41dbe113d1",
      x"8f153978e5b0ab640f98793f03f1a6e0e93cd6bca67e1ebee44d34436519487a",
      x"7b6f9cec34087447f6d50608e05d6a765fe1f4c4291771baf89acb40b827210a",
      x"beeac90c1d5333d6f4b5afc6b20ff032c1c8a03733e850566e53bae4229b1d05",
      x"b5ba2d7d03716ad390a735ec8b8555463bec8b039a7aa7b9752b1957761d7628",
      x"34509e34d522abc22774a4d682fcec793b95efe7685ec81fb9fe6c51cade072c",
      x"49d4ea706f20319fcf575edbccf24058fd30e3592f4fe667cef1ecd7aa0d41ca",
      x"da7b3e8a9168ba6edf550b88c6f9bf2f3db6458a6d52143e97f3c96190c1e137",
      x"8fd4bc0b07220d351c4d403b44feb28a12ec917eda068bbe70f2ed285f1c935a",
      x"ac3316f13850b370e9b64e59e952b8974573430a9c046a3d93598ee67db51cbe",
      x"02e0d0bcc1017b709c9db42fc1b369e5b2bd287486d7a25451d345be2fc4c858",
      x"15bf16ac7c77a82d49b247c9e20fd9f2fdf92c6d558a75077912decbcc2ddc49",
      x"b19f39a6336940ae2e66ce15158fa1d22a30b5500c397bc9b6173531c9679ebe",
      x"6cca291179dd898504862b19e9ceaa61a8943936aa681bebaea2bc252c296251",
      x"fdd2fd0f40f7186608c2f60b8e0ffce3eac98b0c628bd503bf086a9b283d8966",
      x"df38278f06feb7a584e458b6962a57c53d361756243abcbddfa463175b21d99e",
      x"5fe08ce02257fcc87eeb78222da902fa6f3cb5dc92daea040e88376745044bc8",
      x"ef55233df7ea3750cdd9468c94b8e82cc2a004c6bf8aaf19e9184628d9a178fa",
      x"7261d4af4d3bd2d4fd5b97a19d574f535f24b963ba27dc83c3d33e1e7a363882",
      x"a6cda8ac3247b5f8efe9c09ae8ff23de25f94c9676d35ee4c35d0019769d6fea",
      x"7a4d4500d064be781cf2638189f2e76f2dfb3151935eff613e6044a2860f6b3a",
      x"c2a68834978730c6109c0f93fef506528a03d084853ff5c8c7dd6c62f73a3151",
      x"4ef8954f3692ea9e131ac2ad6e9f388ee07c031bbe4c318374218098f8fcb864",
      x"51080de658eb68339d44936d9224798789e4dd12e2b0139a60950284e8b627c1",
      x"b97122355ad8f9ddd09abb1efb95499bfb2fd5cce6d86733427b2ac2f6501949",
      x"73ec6ca28473624f56c460f30155ee134a215bff27f5b58cbcc2b3b6c22d28ea",
      x"9f09cedc7026eac5a4eb54fb7f5f4db4abcc3fca949c3aa255530cee1dfcab06",
      x"4893f86ff189689c853e14931b5e295a498a560c528e449b464b10eb67c77712",
      x"0dae30ccc5dfb2ad5630ffaefad35e804c266d00233d6be7c9ff30fc260bff8a",
      x"c34e058e442510d0bd3f7f0edcfd12b2d11ae479a3e15b6ff0609be10158f0aa",
      x"a073908159740257d408183cd46ac7d7efd418120f5b0e1129ab399c9ed1d69d",
      x"ba49260a33d5a3e98a2ed3ca174c990e7041641a25ad1c860b903ef036ad5f97",
      x"b43f7916dc01ca6866ec94fc909037c4418d5ab24c7b06f2f37761ba783aad4c",
      x"40e8043f927438e1eab077fe4316ae050ea8d45c6e389f65afe763679a580c60",
      x"0ebc16f6cd851f79e89b3cd186ea6f3a7cc749d6a049f11d3a92bf6da90d8a88",
      x"03a5da6243cf083725c428c9b11ac518767e8214527a3584ba33f3e7dfecce01",
      x"38d0e62250ac242e82e4eb2a3b9fcbdf8384b6c268548b2c03dbdfeb22be2fb7",
      x"6b05a1320d1e9765f38e160ca17d4e291e93043c1ec511df6e0863d2f773a239",
      x"c7653b4b6754ebd1bb18d9fa2bbe2827174310b8163b9a3cae8f8136cb3aacd5",
      x"6f9d8a56b73ed5d0e66e5706a4aa7b454fb7202262677e90c9e142fc75a4e030",
      x"8b8e299eda2c1c586a7f1c4d1c31cb2e8dc9e43a966a67467ad34a7c67efdbcb",
      x"53032de2835d945dfacc96b676f6311c39b11de84a0a5e66eb0391707966d6ec",
      x"d451f6b67f33491c143ff3f4317692dd7730967a9098264b51bd030f2882238e",
      x"b49b61824724df70383f4af3eac3cfcfde2fe110bae4e0853ab1518d51cd2fcf",
      x"cb19643c5dd03fca85f69d416650e8109cd071ed7d1efe442e83b7a90bdfe99d",
      x"5e7c42a21245ae788bae00603c547b9a3b82a484a36c8ab150533252ee931ab9",
      x"70cb230906ea61dc59daaeea85288505860cafc7a33083836b05fe229f6823bd",
      x"b56b22e1c72e093d466e4f68de49c22f6ea9238214f9656dd1292f177de09236",
      x"9972fc4c9c65d50b564f539face3ea9d14611632a8177aff8d207d2eab848eb0",
      x"ec3540f9fff74c4093e474e8c0da809b86391d005ab424887dfea4be0ccd6fb6",
      x"a7a4ca1ff902d44876fbc8a4ea71c13a402e971c009dee2840059bdb02f0ab9c",
      x"dd48229afc8e1984f4c92039a74418a11f8d4477910a6a3e9faa99fe55db3630",
      x"620e3c8ca4a97a9fe5292aea06ee4846083f8460432d642f0f63d0b03c7efa17",
      x"b4e9dd23007509e9a151950f9171910b25bc673e732dc5c1a92dc3088eff85b4",
      x"18749a34d84d6fc8b60917371447ed70e1893fe52e7b9de323bbf807fe349a8c",
      x"d89af9ce3fd753598a4507d812a6895cdfe12e754210290461a081120ffdf05f",
      x"e33df546f498b4fe3191c862f85cfe65c364e272eab36af7d4f0d3bf90fee230",
      x"d7ee63fffc3a225e474437ce4f7b8d908d94ee74270091a6571734bc15ff729b",
      x"1cc0418573347daa14de798e32e2c51c5d26608a0ddc6c78423696156db659c0",
      x"ecdd99d0bf206fb39bfcaa288200d99d36af7eff4028c71a98da9a7de939c2cf",
      x"3d18caf5f1800bd72e957c9d0992ab87dd8dd04e71fe0f9360bf313094b0cbc6",
      x"6b1f6bd1bcdb1085c68f2d454e4ea786c2f4a331ab309ebfabdfabd0f451178f",
      x"8d70f29e6a0ebd196a0a3fb8bee9dbc6637a1569d809d2a23416f0948ee8597b",
      x"f4f28d6e91c015954542cbe9cdd2e876788aeed50bbf97d72e15b181fc87acb3",
      x"3bb84f32f4691cb1b100904b9ed2d5ac06f12c10560d0fc55d39e98c00651bfc",
      x"51a04045b72c11d32686183e050ede3cd91b90456d55e61fac3dd514bd0e5afc",
      x"bb83130e23ad32e011635e232f3f75c7866d53856a5e8209fcd98172d687f41a",
      x"046c642176cc81c15d3b6d34d10fda92b62407ac4d81d9f4b57df6b6c985873d",
      x"797200efe45dc0c345201ec70455c899b34c2d41bfaf9b219bc8aabe625a2b1c",
      x"695f17612b27ba57ca4a2ba6f7c75f634eece8f5aa58af17d28ea07dd71e0fe5",
      x"3786ccaa22bb61fce3af1556612b4d150eeb21e424e010db171ffd55ff4c54d1",
      x"f516c61a932203c67fde355768584d987030ec8b550e57a355a1d1518fa580e5",
      x"fab3433416fff69078fc3a32cdd1b2a5d5acc6c717c38d12c69a1c5d008b7739",
      x"c6aa40fdefcaa96a5b76b38714216b5ed715ae3d9f822d8194c4f599b6313003",
      x"23d47975a35453aec65f2334b0e23fee00bace2bbb5698cd29c6bbe6edee3998",
      x"ebfc5c89f1bf309bf7842b3c99038e1da261019eb19d545d1abbacaa2a714cc2",
      x"21fc646c9a36679d2197db46725aa38c3983c03f89d7a9bf04d6ed0c5cfc0a1b",
      x"ed4a977ac42d688402e6ac080568df53fc8c456132c429bc7d4b9c365f7e7cb3",
      x"775b57b009258a10cbe093c2ae3f1932932f0544dec4989b5b7aad73abbee2cc",
      x"0990681981c22f2ae19f11249fd2251618d2835f2cf2c91c3939df744cf30218",
      x"98914af70b423f83278053a84ede91e53ae76fcb7d2e815403dc04c87c09e3ef",
      x"05c2e27f57fb907bba5193323e7db20e283ab1144c0ea9537d48ae0c6ec87908",
      x"b8586156e0d3b18b80289b859892f2a01256b8a4ec608b55fe576265677bee6c",
      x"2e6b869180397be0b230fda724a30cc6c4f01b9a59f5446c608b71938f86e130",
      x"f7d0a8688a898d65ecd16486a1db0d1fdf124eb5d118428bbf6890ac4e4b1277",
      x"e2bfa0962c881263a77a36d02f1e30f7397c3bc13e312d38aa77f5a8a4625911",
      x"5f1bc89653c7f9efe56cd83ed0ce94639f31dbdb225a284ec7a27badba862863",
      x"9cd9b5580ec77518116b7e0720d70724cc980c373171c4e1e50decf298a80b99",
      x"dbb9ccdf9e761ce0338517c862d5ff52908e503bfabffaa71e271ed7e9b72bd6",
      x"249b3b5907085d3c18d2a761a5e7fe6cb476bdeb440ab4434a39623ed6ef6d83",
      x"f703193881d6c3953634a624aaa5b826049b4eb83f7e771865b60c3c3760ed1d",
      x"67683c385c3d514c0408c0a93f3f26c5542581c6c04a9777e8fe34f7345ef756",
      x"a0e8d442fe5d8f59e75915e6ce5fc8ce94bdf9023818f8b970a839c77c941291",
      x"e490ecdf3715a512d23fbb8184808cf0edceb035593cf103d047139039dcaa2e",
      x"ad65e26c485e957ebaef32a93c5e4af4f720b2ac46f5cd4a06375baf05f77e43",
      x"2d541311d31f4c2badb7c0c98dc268e5795ca6c491f5f409784e52aeed37b98f",
      x"fab5a9dc7dfca9df353f72447e975526aa8f5bbf95fb70b8899736ef5d9fc29d",
      x"d2a6dfa2ed57aca0a5b48eef0e4bc02f3f2a3a72c0bd51229f401a5ab97fc424",
      x"6c37c608131d7a7ab5443193ab45e15db12babf6052c32144a7a607cc0ea5a90",
      x"a7311054b87ec1132f5558ecc3626b3026f5d47418bd24375cd793e3842c2139",
      x"6d24770e13639e6b84c9b87eeee88f00418f39bb1ec879d9c64d39c76d99641f",
      x"acae870721bf419d0bad092c73988ffd4a1ae6e3ce22c10063f19f309fd4ba9f",
      x"9952e09995327390d2a08fbb2b8fa95a91c3d257fb11dc617161a2e33faeef42",
      x"8a4bcd684690d2f80ee318164704bea76fc5b9e1689724830a6348c4281c020d",
      x"c09f5bcdc4d330d24ad942575cc15679c7701d649675cb3ea786015686711e4c",
      x"ea527861b97403bfcea694ca12a749c26849af363b41d9c752ba19b396cd3eb2",
      x"bce303b729e4f4aa57f2d7349a71b2668da5c21dd4b2689d43b5c9ab72b23a99",
      x"e283ad0c1e20fc03bfb6050dd8991e1c9500b3157f3885e88699361d2d08ba80",
      x"d45b2a508fed4614029994325e7cf4ff97b79677eaedae53001f0ec0af024626",
      x"e66dee7ada33e1ca287f7f0d6df70de42f9fbec8933f1bf7376f5111263144c4",
      x"ff64930a5f67635077ade2105476a62de1756fec374aba55569019180080d09d",
      x"f4a94aa75bdc266b19d7ef16a3f4fff2f466e70e054c9ee003b9a7d84de5b6d5",
      x"265b6450a83b21d46d3515b17e0da025e166815d69afbbd72f47e7bab915b691",
      x"a35f5fb09c90d5569b37ed0d4ebd0067071a2b3f53e17e37ca23883281003ba7",
      x"9b4ba956d5f8ca0029758ba492e4e2d2f7c22f29517b93f59a15451bf3f78b0b",
      x"07d0e210cb596041ab311b461b32934c894a453685b1c358eb9a40b57e0bf550",
      x"3e472c4a760c65240b5e9e9b4004bac975045505994f01fd6de78a04e78df1d4",
      x"38e2ff0fa1486323a19f08a6f36e666fa4d0a0f07411c4179e3619ffd6aaa4df",
      x"72f6391006df2a3c06e49ad413edfe2cac18b02af0d4a050cf74d842960e7197",
      x"fa9d742b1f09bc2833a1f6afc68fd6c5bb5573de018335c79220a778d4766a61",
      x"be23b9c9fef1d2f67b416c49bba9322c6cf131cf498bcca718537f2fe91df4c1",
      x"d1c309f4dd3fb837af4a8a54d942399fcd82e6eae57369e38edc7bffd2e72718",
      x"a0a1356613105c5ca6f91d69f6058060ba7c77cf1c1b5b565242ec1257b68f3d",
      x"fe28472936d2881b04e60c79fc9dc85a8fa9de2a6ad5affdaac26126bc8b896c",
      x"d9f7d4c60e9221c50eedb5ec5fb886fdec014234a07c9e59f319ca655234655b",
      x"1977164f851e005dff3a64f9033faff5c3c6b77530461c7f2e20aeebfd67ab22",
      x"0f4ca47a88acbd9c5d85fd6af545bc5b1f996f091f71fdaa0969b2df4a2c361b",
      x"50b8aab98511f7edb2ba5ab8fc9d7396e9869ab11296697a206ceebd79aabfa4",
      x"849a2d5edcb3b3c61aec5a1c9cbbe7af336126b287398af743a45566b0d4160b",
      x"d19e7f8f749b16b8bb54f5d3fd954cc163669e6fa84e056feb235e212d47f3da",
      x"208c9d0da7116cb38c23cc2a70abd5c757645787e9d23175e2340e68a543a8c2",
      x"690a54f68290df5caa38d1aa820ed581037e803c0c21f7ca54e34493e0fe1dc3",
      x"50c507faafd402e32125d97dd973fb364bb59b325aa1e06f6d07a3a8a14185b6",
      x"8f6d9ab18bc4d9e0df447c39cc6a4aec6f37a747a469fd492c07fd2ad3c58156",
      x"b066d506203f8d947f968f1dc844aff4a3e32f802430ee8a9017a69dd79acd0b",
      x"fb69734a4a24b0d57eb5244040a1e5238a12917edb0ef44dba2dfda70f7be842",
      x"4d8c37cb9a347d7f249e2e648efb565eaa7eec635160c41ef888009082a07e11",
      x"1cfdc3a79ea4d8a31b7173332cd7a02b140abbdb93c8c66f51b4f2b48642e066",
      x"7ddb1c152043367e45c23146cacb43d8741ca3be49eec7af55988e61b26c14aa",
      x"66f90d76c70e73700b728f5706877b9118e506003cb0dbb17c81f8d916279387",
      x"b0a05eff22c5f6a8042f5c2807a54a579dfceb8713cda62479c7be9879970116",
      x"3d6252ec7a1dacd6d716e8b77d65be17e7a3c0fec089a9f976f3d3746c471780",
      x"5371e999012112af25a6b259bfa234a194de7a56a477e518ebcf7ffd07bf9dd4",
      x"2b9d989d98ce44dfecbe525a504975ca37f74461bdb7d243496ebf03b4456e99",
      x"7f5f01471c595cd46c2e5d7cef35c62e8f1b391745695201cce65824d7324245",
      x"0b4666fe8fe5afcb259afa876113096e42d21c3300374595c88a54ff8fe54c40",
      x"2a6e9e5b3620ae434886fbe1a0b768c02981d8408f3c1d49790fada81ba5015e",
      x"f029b6bd25241bf5eba358f803d37acf00e87ec07d9225330b5a6c06aa29dfea",
      x"e114a9d3c734a7c135d65f917c9ca3134af8f76f2c390ceac12e4594a039b462",
      x"3f164f3f119549ee5be5d9cc317718859ea18246d8958791f092a8d47de43d04",
      x"d577b3a389a3e80de81d702b5e9c45af454986eacde6714eadfb2d800bbb9cca",
      x"30f5744590382942d62107e9f6e9d23059e37c277a42d245e58864c6b2dd53eb",
      x"d9beaec81e1a3ed12978a99d3a8027bb2488a71c4c195ff387d21c43203b89a6",
      x"3620085dfc7355f61e9169bd7275f570631f579bd19ee456f3d8dc6dc756d61d",
      x"bd93b31242693e946a6d4ef48fd89d9ab7c932e955ebcd74ab508df89c171a6f",
      x"8f349f93c3edfb5eda3ea9397839663fdc71bd052653fc25bb784107b31c596e",
      x"8308f79806ef71de05fe7c890726c21a93ccb99627ccd18ba408d462732e9e51",
      x"4d60aca89fb79c6c0d37cb5fc8cc305debcef9ba07272b88de84f1669227c8d2",
      x"08cfb215c4dfec0154b98eff71be6663a0490b586036ce898165516b3f4de157",
      x"ede40ddf01f2105649ac5600734ed31f4003f3913d44290144dc7077dd0bb2e4",
      x"6e95d5c72fac85fd6650b7eb389ff84006625231a046d50603e0ff9c8f3aa6f1",
      x"d34a0252bc902a3779d9db72eb622f7c80d744dd0702ff8f5b3c8d254f7646d2",
      x"4bf90ff2da773efff867cce12171748e911fa2438ad3bfd20125c0dbfcb93f5e",
      x"cdfc13fc9af721a14d933d82525d3951842191d035c3929909cc390c1b40af19",
      x"e64144dcb136226d5f3878d9c112db0ba9cbeebb804e3638ba06685cb348fc6d",
      x"d87b27fedc8ccd8e381383b4ce220ea2fc6534bf89a1c624288362d9c318d636",
      x"c059ffb0ce8063fb030311ea991a259d89a3c77a997b4a6ee0898553285b45e3",
      x"66b1026c21c73de8d3d362fcb9247e9192ba31044233d3ab4199ff1c622131d4",
      x"5a70efc7f35fca9c574be2d6a8a690ed58529f3031fe7f29655cdbc9cfbf1096",
      x"db7e0a8ac6788e8cdc966b9806ed55f6b4b78d4c9f6ccc466fdb5facf54f6f92",
      x"29d484ee0c4d6ee1411089eedff481ddb2679663b83c670ad3aa8101b75a575c",
      x"44d2e5baa5c2d42aded7525e64ff6aa007e4414e37f283bb2c060eecc513a17b",
      x"b42fe3986942359e4b406aaae0882874c8f826ded1275dbc496249dfbcafd212",
      x"822a52dfd0f496fd5ec4f297e815d3859ab5a2c36672f990af41f3eda346c342",
      x"5ce4b1efd420525a746be9b6b842cef0f03c3bf5a999b3b27f7259c2e6c2dacc",
      x"1390b3dc1020573e5130c8e8c04dc85362513f84a4982a5c768adf5ae28e4190",
      x"0ee0489a81b6ca0ba1a5cbdbad7245d534879bef3338d0703a0521662be9bc3f",
      x"ccf594ec8daeda80f9940c83fc89aba90d7132fd12243598918b3d91eeeb13a2",
      x"204e878e1649724521513daca05d8036126c90304d030e8c7f4d79c0382143dd",
      x"a5821ffebc7e167ef8d34f7a25ba13412c9ce56c6ea297662e136c77a5dcc0e7",
      x"5d2e703b3cb01d8048aa9c34af639a3780b18e4da5b2c0927937e805f5b60ac8",
      x"b7abdb522949e372809dcd4847022619dac230dde38aa235db92b927e79d4f30",
      x"75dc05614f629e74db17d7f9821bde59df5edc5a5afb92bb783bcb18d1e5089c",
      x"4c64a9f456812133585ce359dfacb914a0c908d2b90b8dd28086236bb0dd2bb6",
      x"14033c1a4a42b18f9ef18794375bd3530a68f53b97277385c1ddd905bc8ec3d9",
      x"b29c06d49c941377bb5247aff0883419f394ff944d140e5c04f57abc51db0f9d",
      x"e902f60e6fa65ea8a5fd2499191102e13a02a3e5fb95b1cc174ab5e428921703",
      x"4d55089df92035b6d8446661864b72e4d8cad4a384c01ba3f6ca285eaea9d293",
      x"347455ff65e80671e7d2a54a30bdbaa388e99d44766731d7381ae91272e44e23",
      x"1e75b068e69d7f78972d6ee2532a100120895777a1c7fac83fb24e24c278a055",
      x"5b6e8c00c1f4090f59d9003e78a0657443eb102c26a6136bdffa6ad55f098759",
      x"00574ceb800704e6123646384fc0eba88073039151c2e96b4751b996d97bfc1d",
      x"0051182d8875a88ecc0fcf4167c81d01e8324256717722f82a7b61e5c6a52151",
      x"e8f46a16a083ca5c619201b38b0ec94c0cbe3055afb1f5b15e3902e6c280ba1e",
      x"7776f2d9d12134ed40057cb0fec599d869d7f3d04d5bb09e6c8101993e65fdc1",
      x"e3a9174587ca23729971492af8958ac1ef011e0cc9c1e5dc9338f46a5b59b7e3",
      x"5e08812b4b4376848179adea46c0dc82494fcb18a6f31a4c5177d3c7bbc2cc9f",
      x"1517147d05ca1479213e49143f673efac5ba92177b05a16cee26a17557f536dd",
      x"060c3a9312091abd94baad63c2124ca0bc832c2e4486371b6af436142d21b34b",
      x"9ab6c8531b97d0a4fcbfdf613b50726dc03f665507f9bd5ce4b1078553ec37af",
      x"9cf352429281b22f80e31b088bb00677eb4baaf61392286779bd579f7105d6f2",
      x"43ed95fb68ccbd5da542a8a1f2fca0e41c346707ec9c3d22de7b61579c573ac3",
      x"684942b362775fc9af95be14d1abe51b31e0b1106ba94955807c4a2856d0c5e5",
      x"50eb08f403227ef49b9e339ba4b2e1b1bbf792f35224059548a95c6390fe048a",
      x"2799f3d3da370b425b81b030d1123fdef61bad5de9505df6ce8f3a5c3da6ebc6",
      x"7bb0e2ed601fbff6bc06cae1a9a54b34faeb63ca4fdf06625f38400f58186008",
      x"7af1552d07eaa3d516747767f1ad98f6793c12bedeaee3b0b0043b3a3512198d",
      x"465a7a7c3615fc5acbe3041cf441975ed04c63e2dfad09d5c7b12746507b252d",
      x"4e804dead732db638bebea85dcee35e96c15702e268924873b4b8647cdc4e7cf",
      x"17eabbba1bef46a3a87eb9726168229115ff6a5570956ae911e08899d1c67f03",
      x"b206c9e20ebd8f2c0d8440e6412d7190694fca43cb84e838278bc0af8df08c49",
      x"dd34a77c9b5e8a62639042d097ffc78dfb308174f03a4d3a52ba4340ccf39fa4",
      x"ece3da863d4c90d73b6171423e1e698d9888d852f0d95018ab788dc2aa5fbad6",
      x"65c56b213f18795b428e45aefd7735dff0e410236e6b09f8e4ee8ec1854c7e43",
      x"cf2d87f724eb29022c16ace76b66110d1bff39cf485dfa0ef09f72462787a744",
      x"ae8f04e35cfa9a8d3a1856b37276607a7e690ab9a359ffec0d0d29e36c486e65",
      x"e9a35a11aa5f48e024b52047de079b66d41fbfbf1f747806eda41f19e1c629d2",
      x"db22c4371178687ebe4e1f8fd34c26110ab9bc18f921c230623f9f63e6809b41",
      x"658861aaa7ed6f045fc5940ca35fe95943d06f44d538e46c3196515bf823daf4",
      x"8fd0965f955f3718c09bf3797e2107a5af4cf3b02c3211f05ed4cba804f66948",
      x"0802be32d57178299a518aa2ef7d716ac0c7e0072bb9acdd49123b8d392173ac",
      x"7bf7bacdbadba7f02e6a7758ba8f18713ca9a9c8a6bfabe48dc76f101296690b",
      x"f23533816f0bb0f90b7c55f39ca96de07b9e64eb70c0cf9683068c90ef59c3c0",
      x"b695499a632ad7ded886ffaac387963454f9f7a27503020728f03dede90ba684",
      x"8eec3e5f3d309c24de0c4fea1c877a27f48f2316573e85637fd6e75db931a736",
      x"74b7a8297ad10976fe3cf81222066af0a911e10c3c5f488e7fe81788c9c7d924",
      x"d4a3c41f6eb5d82d27c11af314bd1a4ac895d19fda8e0c7889a344790d7ad43f",
      x"65976a3c34de4bda2ffa9e7e5e977f649fff2daa2bbe8adb1c7841c06d0a3c77",
      x"7dcf0086625440b1324f1b98c4d037189c5a7c27c1ceb5c3631d9fd51364c26f"
    ),
    (
      x"82d6814aad45736b94325e2a14a4d713303ef4399a57189606ac1f4d0d344790",
      x"cb3574c0c0aaa25b3eea1a4643e7d4c9cbd565119c6a546f43bee029b60f4fcd",
      x"ad2860b7576c134a115e7c7bc8b0dc6eb49d0a35c69f187472f3a4065ab9a5c7",
      x"2ba0292ccf909c3017c9f77b78c7887a2e0b56d700f99d8e0574726ee7036f1d",
      x"85aba9913bc045add2dd8e9e638e38ab6f10b03588179bb06086665408c69c7d",
      x"a30360192e6b3983bbd73fbd710dd8c4da8576e42d06bc8262ce3a18fab95b11",
      x"57df892381c90ffe7522a03248ff9868e4127a5e8de5394a5c3f5d8c164e2eb1",
      x"45bc26911a08dcbbf7e8db4686e8b80c68c53e759b09a2391d68f6ef7aadaacb",
      x"886939dac426a389d69f8b841ade3c79e6b1254ae7d15e789363009b16239c36",
      x"e30be5cb39f58c10be7fefbe5f52e0d862686e8bc3aef09e55816eab5a8447fb",
      x"7d732c778beed7465f3c874f1ed5884f1823836c24a49f62d19f63e06763affb",
      x"3789dd427c29b4a49c12a956546b5585371ea6257e5477d0964c24e0fc3cde51",
      x"640c1b9867c1e06e216763ee8994d12a8625b5b3440d0239cc4e74837392866f",
      x"b3acb2d49c831d1aefe83789df965b3899af3f7ac10252a175a5ed5fa54ac2db",
      x"dddcdbb5a308c061c932bf4a36d262c6c74eb099ef7dcd1d70054cef40ef7fc0",
      x"289daefb2be87da9dd627f7a781844af3ed83ee3438a775e3f75d79c69f68c87",
      x"8480c531288c180bf6de38411c1e8c884f7f07520894577b87616d4ed942b148",
      x"f95509393addfdb61f1155503b50c02bbed6c678bd9169c11185106f19bcaf61",
      x"7cc9c4c9697605e7104015d61b955c3b2cb7ba443a1da343228781576cd56f26",
      x"d282f7cb5af7206aaa817a30f5246dd2d4427e75d787117b42b38ff73534980f",
      x"b6587ca4f5e5bdf444fce4ced15958ba79cb537d08dced35ffc0d3d1991a8e5b",
      x"029dbb897373c38c38577c7a2c68d8c6f0bb27534c3a70fdf1a8aac9d344d883",
      x"e65405a055b60ce109b17b491912fe8ffae42ef8ec68cb8c9e764f43dcab3e79",
      x"0464f4d07d4f60a05c0a2cf0b82588507db49dec25c76f14ea5ceeba8914044f",
      x"43d97957745a1878ea6a0cfc1558017518af2b5e3311529068a8e00eda45971d",
      x"18835a469b1cad89298295b59d7edc6d16484f58f2306554f25f1bcb29428f2c",
      x"cc6abb470d67a1a38175f95eef8d1281a34df14b74e453f7b61583bc0451f526",
      x"3bdf31a8acf06e96bffe27c2e7ebbc04a48871e4ef581cb98aa646cd11a9d171",
      x"91e8d531ab70f9752c7af68703a4a3b3c70bd5ae521d421eff1dbbc86a91439b",
      x"c8912d793b374c9576969fec4a1f27152e2716a24135848b1bede785e44dfb1e",
      x"c25d56b164a1d208b7ceaa72038b01a87b83a8abe02fb8772fd6af2038b523c3",
      x"4661abafbdcdae2af852e432957f981614b19a9de382d0fb334ff18e0b0ceef3",
      x"7f840c185e72e2966bebbf90df81568a4bc5b4c905270af945a2bacffdded00b",
      x"62378431f2c838684c83357cb930fcc9a670dfea3ebb9f5b1d3a70c1a1a78caf",
      x"81df1dd291c7dda281b95dea9925f990ae74bc2095f9329724ae5bf688dd5d9d",
      x"685cc6b4d3d58b5445e2770078f33d483a6429cb27db293bdfa69ef71b4e52cd",
      x"e209deb91a1e29ae6523bc7509d8fde7687cd3145ad609a4e795a88555684c0c",
      x"d877c4717ad019948bd1d4f1b8cb22f02a16814ee3bd426323c11efc67e52592",
      x"7697446540950de26829a949829ab90a3f55d69d833bc0d5baa80c55a4f08c60",
      x"01a140cb0be310f777d0a05eff44bddf5179259a4a8f76a779dfd5c999cbe01f",
      x"53cc35d2ab81cd6e6bc00692e4ed877d09e8ff9b3192d84a705cb97103b12bf7",
      x"78ca68566b4fc47274765c5dacaafb34fb7842e08de30874265b15dbe3b1a79a",
      x"a7bfd5e1776bfc926120210c2699d09034552fb84eb63627c606ec65c812025d",
      x"ad43ecc308ea0e5da16feb713b2a99b9b1af1d3ed37bc69e3502ec54af2e87f9",
      x"eab3a1a05784bcc23c9886d2be96a7c8f6355545fd88a9d9c0a6d68a0174c657",
      x"040a9468991eac2e63657b9d5c4e6a3d3d7a5075a1f6abe4c0e3367ac0d3768b",
      x"47e98b784012cff4943de760e789c3e78d4244c36277fec513ddff311c411f42",
      x"5a66b5d665c160fced4ffc707ceeac068b1cf40faee680730b7d5ace7c04438a",
      x"808a3142d10888fd750e6c5abab5074021fc7c64d1d3e9800e8bb48afc97d528",
      x"fb78aba4d20925bca0cef6bf1f84daa460dbdb31d38d7b69a72712e254c11e0a",
      x"4a04a5b6690bab77b07115989e9e7090965ac5acb6957d335f11c462aeaea295",
      x"e633e0618ff54d1f944a97e5ade1c8119ad6eafd1c5b761f12fdda65d8143d55",
      x"698e584fab498693959dec7d1842ce8fcf15b3316f6374629c070a64ecab7c17",
      x"f0cefe6b1bca1e59b10a8dea2f2099e595849dcb6feb1f250b740b77f7b5c624",
      x"cf67c7bf5572e5c42bc1edde4ab43b7f718934a7b28ebb5832e74652e15d0534",
      x"1d87a5706d9e3528afd5a8b1656c250ced26d180c6d3f54f26905a81d7300e6f",
      x"3ea192db51d2ea5abb698155ea239cf14cd6fdfcb5c104e2ef3a2b20db1cb2f6",
      x"870757b67ce15d26f7d07aa55e67af822c5e328c143004ae5cb998b448ab80b5",
      x"6e530dd57275ad9acef579a48c40e9dc8699b26339e77d7adb2e947896251ca4",
      x"b461c11096a5fabcaee1871f371de7fe95a66dc4e6635013930cc5935eccc0cd",
      x"ea0627a6c37de5705a062b14d6b9ab88309557c6f43fd265b0088ba15c44ead3",
      x"7285cfa8112b7bf9196d578b7cbe3a985ead0bb4076ece43a4d3f580fa1b7856",
      x"f2fa7c7102d2368b47da571a90c42d29359b683fc450764fb875856e5f2cc494",
      x"04a5899ea656bc2f97f51f0502a537e4a77e516601e0958fc7d2b696d2f71c30",
      x"7ee63bfca5a4b9b8d96271009b24c325d4b4c744dcd262f1c116799edebf00ce",
      x"33692585f4bed27117a33b9dc1136b6c1f335d3657b34b51b839d244294db248",
      x"7c9c3f8056a23cb993aff6d0cfda1cf49dc99d366a701f078f6f29e5dcc0023e",
      x"fcfc4d861c858f42f2a1fc3fc16fd4b189371408aaa171bc6cbbf262b29b91d7",
      x"1c4c650adc5e40dd890ea97f6ade2c6705139cff9a061573d7f90b7de3a3822e",
      x"dbc10696e7948a06c031a53e3fc99ce15b7b692ddcf169a51c871ae493247752",
      x"cea1adcd6442bae22f23d8100cdbf1549008567dc6085f4faa5672eb68383cee",
      x"dab043223148e8811d9301e5559e726158d1cb58a5f8994f354a6ce2ce1ba7e6",
      x"ff3f9c49621dcd3efe45a11f5396629b7aed5f39ee023a3d7f71849ea03c0f68",
      x"8a024666256398d5ce6f0cc5b5d23d31af2e875d29519ffb15ec27a094dd58e9",
      x"1bc88764d6bf41e2a3a18fc2dc6c2be4c206dcb6fbbfa5088e60f8ee4f50c5f1",
      x"e41e07c3587d6e8dbff3b66f97ce7bc8e2ac5b45caee1d2402e495ffa780e5e3",
      x"546d2a523a3a711b0908e8b950a9e87ac452e7b8105d06abd14948cbdafe9f58",
      x"32b9e321728935b86cf45522b673cc698e31e6dd4ff5420f45c62b4db1453c59",
      x"a79b90a0d5be4def3d29afd69d7fd4cd25f9f4db7abea5a758569defe52ab4da",
      x"2d932ce09ea9ed84c07943557d94f87221829058fd8b39b6d575e0785f7a23b9",
      x"04be0d0b8ac89554efd1e6c4a4a12908e2226881e64dd613166f9189289a6fd9",
      x"92ad42b9369e7926023dc1ad8e0932cc1e6f14d4766b00347a1c9ec0aac1b258",
      x"8a8739b84d467d61179eb88a68cc5a86f6b6af04a35d35605b03e28ccc0bb483",
      x"fe0661700db442cd79ba20aea02c24b7ed5ecd7f51c53edd1dd2ec732a265541",
      x"4c332268487574da85558046c4411c4c6022183e3121c5caa9f1c126609390b9",
      x"82ef190f2edde0afd3ab4f6f627a30dbb1fa2da5bb88ee74cd1a99dea2a39dfd",
      x"468df61cc94cd8f434399c15f35bb52aa5e111788e9eddede2b7dfbfcf3345c4",
      x"87b27d9304ea50a199144ab3d5565a856446a36764c7f7213df435c266ee0440",
      x"3b056f91d3eae2f038a1991fc53fb5a138147d14b88a473cb13e120ee51d4e6d",
      x"c5fc1fad5e642fd08cdaa36d6012451100daf066981bda7f0f46b29dcddb5262",
      x"37a5adb0739f5aa0834f67ea5747f80199175fff380587b1bff162aa59e9688e",
      x"de9a8f9b887b1313bef3189bbc68ba1abb77eeca185f4d05bee9ea9cd215d1ee",
      x"4298ca9f129d1727208aca82fef6cd1ec67e4d12cf89c5b2dadf2e871463c2c9",
      x"c7e79190aba12ecb9ae198fca72cc3641b238dea3cacfd71fa065cdb03c39e61",
      x"61dc58a324950e37870c8b0f3165926ac9037148f951eae4a3cb808574a076d1",
      x"4572b96486fbe249154dc0a423564fec1e662dbf47976ef0abc27d1f22f1429a",
      x"9a0c510435ed721d0514bdd582bbe23fe2af04f62873496fd7d5d09ef3cc0af6",
      x"31187af282980d65a66e83cbac71d4c87630fc66714e90392465e989cb29254d",
      x"1a4f109c8c6d4a304d6198ebe1d7af397b4fd84b20e9970c0627746557152fe8",
      x"f288882bc4498562691ce39bd50ddcb5432f9d6f8e9a43f2119d41ed874d352c",
      x"fc449751d87dbd16d9c3ef22a598a9ad584ed916d3be8701b424236d1fd85211",
      x"0df24e8eab1ee3c4889dc30549887d14397e73d99c125cd81873d46b7a59d017",
      x"6049caba54f32ba7309620305cedd9af5222e64c98255d30d7ea2d7b8bd0da0f",
      x"a0518907e881ce4cc61614c9ab06bd72f4a3a82b48689c05545e3e8c1d1c09ec",
      x"b58c032ff0f5f40dd35a1ac5b033b39be531377388e3b4b4b00ecefb443f13c8",
      x"15f2af212f4e93e68947e31ba30e786841ec2adfc65157923d56eba1ebc0c679",
      x"fd87a2d9393588351942bc10c074c4303651644053f58a0ba72a0dae3a9eae65",
      x"eddcf5d2b4c4f21b04c58a024b86d5c47c6c59801cd3f3811b092feb6b3be19d",
      x"72b80ffba41d2a84ac278aa79697d87f1d990cd94157eaa0007f4efde19af105",
      x"630a9c9e13e145feda9bf37c253ca360dd6f44984f4472b01936b51ecfb8f960",
      x"c0be7ddd8e54f85743d907d3eff47c02193565334b0500c66831d548d2539a47",
      x"2d8d53cbe3daa7d46d14f5eae9a4a9f943c7a72eaa1d6e620de7193650c33f80",
      x"ac8a6b49256c33c1fb063c3b2656138b0028d6519caa15ca9b34b8b10972328b",
      x"33bf0a3ff49c70db662a6a164d45a71f73fad7dcdaae16b4973553f7b93ff1cf",
      x"69decce27155eece39a2d84b3281a1ccaea8f93576f94314645580a2db86ac2a",
      x"2c848b6b1810aa97c91c0c09d967b9852acbd998215870dddd7d582ec1f9bab3",
      x"f074e411e2fc8c5a3dfad6c8067a215e8c884c47d357a5e3218ad058c807bc64",
      x"6d31d39535e968274cd4f8b59505dfa1a5e723208b32d3916b15b292e395ad3a",
      x"55961203838800552cdc3ad0a56647af20e4869038637eb6d56daac0c4202e0f",
      x"1f707d7527f48c2b35cbb620450c3568d60afdcaddedc703f25fffdda790436e",
      x"5255496253c723782f96912d0c29f7f4c339fea1875b70913f1b36e4f1d7f719",
      x"a9014e8baa347f34c6133ffeb65c0fc2cd61ae0845c46c8aa488c5e94401c79b",
      x"0e85a2cae42ec87592de62d9c42f805955dd8d423ca66bf903531104130aeb71",
      x"707317c3d17eed73e2203fe06035464f342ede847f71a55aa4c4f841739a12b5",
      x"2371bdd81143fb5b2f57fb917f843236066b93a780dc2031c2d20cb5f0343eac",
      x"1da2a5e6908de506025b5d977776f5fdccdb282cb49c52ea752a4a299617f161",
      x"3decbd4e3a49e604443638b5d4357d01756027cdec415c46f5222800999072bb",
      x"c20bec081aaf0eb16c93ff61c70c1017a02f771d6f7f2a7074e83f1231a6c23b",
      x"ba06c5b44825dc14e8f06d1be2a476c138a9f840e10abc5a6e4ac5765a700cf2",
      x"bc4bad9922b96cffbd06e09f1ce9951cf9e5400f7245f16cab8de0fcd175ef09",
      x"547b407dc71dacfce8379cb24e69d4039926e93c083caa87fe08a4f2b29c07c4",
      x"26be833d4735c066b3e39ea77c4c3dc278cfcbc91b90af5a47d315b6117e9516",
      x"7c91a3388e40bbb8936ecf9d4fe0e045317337ec5fdc1c794da6cc7b8d67502f",
      x"acf991648177f4208cbe799782fd7122f088c8dd204994c4c9572aa32989148d",
      x"ae116fcbbdfbf3b878368b520a0633d1e236ef4102e0a61849ee48d00679623b",
      x"f2e1f7f0d19407755d9e93bbb15f5ae6b70d0af86da3a778cfa301ffbce99deb",
      x"d7965661e46e4425f265dcba2fe839b1aea32816b8729f443fb100585d09c549",
      x"d27a172af546c8ca2407671bb6eb103abe94dadfc69edece7ff43c3da5f8508f",
      x"21dbabb71e603e49133d141ab14be103640464ff24f62d2e0de04eda6e413117",
      x"50b2cafb9a08f7aea984aebf5f89cdf06fd96675b5038149c91457c1d3659b62",
      x"513d63157b51fbb252a42ac469bbebd1536809c33bdaa854177d4d654f68ddaa",
      x"35aa5a39873f9eb5043e0391aa8e9dcdd8c0a37b6e79992ba6641d8cb3cf7433",
      x"d73e2186ab0949392ce88db60f54418593ff4db22ff11d7eb953b72d88ee2719",
      x"190413f41dd5527f1a28dc3788b2d65a625c63afd4edc1d0f979a151e107f257",
      x"eeae413c65663b3bffdf6cc2f7f576ba05f961d8dfb0b8cadb9a16ffa441ab82",
      x"ced1cbcd715898301bddf9349708181ad2cb48a3540a38d45c4dafc9bcff3dfd",
      x"91fb26ea19a93b1f6ebe3e39d0734cc563fc7664762692ae89695b64731d23c1",
      x"3328540a6d1bc95f6f03b5ff4241a26776ddfe688d210433b46cf8aa3e4a5682",
      x"7c39dbfb54c878d60049d5752ed31df92e501d6bb158a39ff4eb979bdb2e1eda",
      x"6e10544d4e744dbb1aea5f274106dddd49def2146f1ee3566f398fc1018363ac",
      x"dffe356e6ca23c2890f76d5801ae541fdf1de52bad19f4d5d658eaa455d237fc",
      x"d5c4fe0343a1e5c03506433073c8c2a59dcf5a628df252348fcfaaefde56e3c7",
      x"e1b3bd7664c04f39f11a04081b6effd1ed6182b5b4c612165f75f195a63cd7fc",
      x"49958e5075e3b5b27375dc2500f3baab0a833b9c50b979dbbaf5b3136dcc6993",
      x"4ffe1245a87271c9e8606f6aa5d63dc97b8879c733fa25719b02fb399a51ab40",
      x"0a49cc6fd611e7b3b70f67e52520f70e3c2f5796ef4f0ffae072d215450d1d80",
      x"27aa1ba1b98b2c9ad0e664955678d0d335142d81f24b69496e444466a510cd88",
      x"b1375b627e8bb9c4b0e3b4d9df5fcd0222059330421a1f7eab8fe3273560d7d0",
      x"35dd4046b35d0017d434f938ab16a57d8950d2ddb0f0e1d9efcdac6c1625e3a2",
      x"13d513f8a4aeb1facac0de36f28d0efb90ab6c8699026256c0eff20fe16aca89",
      x"3ea5391ee307523a868a93ebbed26ed3d49c302c9498891c85dae0a5597938ac",
      x"0eae7ed1af27c8265cde5ed7ac3b1038fb7cc66f171ed7a87ffa89e5a5b1cdeb",
      x"385730066164e5453fd07ce5993dc391f88d311061335e3d247cf3f94fc0526e",
      x"e4f37c291786d446f9b98dcbf827e003e308225e3a77f0ecdcf74808d6e99d69",
      x"a67c4c9f477c4d48a3c34ffd454b1091779b8731143f202ef7014687dbc9c4f1",
      x"f40a2c7631fd33beb49dbbc4f4894baf1aed49e021d3991fe5b8922a10bcba90",
      x"a6777c5b5043a683508192ba3822bc4e780745a0d73fed1b97914a1af068c898",
      x"5a7cf59c334abb1dd4f353685f5483c1d08b56d83ede831c3c2b77178b4395ff",
      x"af08b991303fff41d6ff00379c8bd1250985c349dafc0fb6b2942f3eaa0d8e9d",
      x"39ff8eb442559a432bd29d78dd7a2596d0575ed61e5ee10251517fdb61bcd37a",
      x"f502e2604c6266bfff3cac327bf30b4634efe3e9575d3d21c1f7117019a218a9",
      x"34da324fbf5826d24e845f2e4fcfc4c2047f76116d5c86842288593cbe267678",
      x"53b36fb1ec9a4b5405d6f7b9453f933324a00077cf6160511187403012ca37f7",
      x"4c27612271859c36ec1e45138c1ca1b3c4916dc9880277a49f3d5ffd727b88ef",
      x"d864edb7138393b6254dc1ce8ad49c5be0926d0a317c1e41d99cc69869f248f4",
      x"6d555a94e95771c7c0c173e95ba1aa7ceba1ac5c2f43ac2a5da62623647b67e1",
      x"f6dc06d86c91ae70d5f26bd525dfc6c70fff0f2a87aa71fcd4354a785cf884d3",
      x"fc99a24af4de31864e1ba53b16f3ca1e1ce92cf86c0971dee8f5ff74356e9d3e",
      x"0ab1a63114588a918c00bcdac991c8568c2d14f38b93d5d3dd21af6bc690f171",
      x"233b1c9c94f32d938035bbdb3eab31c07750fa6effcbb25222beb66a400347b1",
      x"c90bf947ffb493bf725428336f79434e74c38b8f54bada5d3002062fd8a2cc5f",
      x"0e98e5b0e9348c577b17112ae75f93279c34f1bf49066748dc4b9d85bcdc00c5",
      x"5384c33620775cdfe5fc5643e6a7cb207253749ffe71c41439ecc5d7038f05c7",
      x"7183932487b967269247f832110938498811f869f1328fa9ad9981c76a9ba69f",
      x"85e2179f46d6f2c3bbcae679ce401978692aa1b867de88d32990a3d2e0e25f4c",
      x"deb3a1c73aa2383530416d87a7b1b1afd87b91df4a661289a65d55b96427405f",
      x"bf4a1c4e450fdbb220a27bd2266639ae25a0f4db507e9241c5e0d3c388bca29c",
      x"235283e808e47a706764b3233096bf342980e4cbb3412d03427ade6091003f15",
      x"4d9adbcf22d5950055aa9c6be0d63851402df1f3b8fb420966dde4bcec584074",
      x"c0d37c93382c5074f9f89a929a58c21a51c0ad61a2807a56057b68918d3c0eb8",
      x"33bcab5c27aae9b42a2c073e994b54c0204cc9a20af10bb336f35fccd999f71c",
      x"8bea418ba4d4b5f351d86fa6d05dc286f29698402b8c156151c0b23679d44a99",
      x"42a38f0b998e691d0110e594e7fb405b64c73002476096ee7e78dd9d69b594dd",
      x"16d3617580fbd5ab57da9be993bb6bc0f93150d02688db404f18fd884f79ff9d",
      x"00782e5e99fedb56ea26925e9fbe3839b7e008c8f40468aa6df3954d7b652e0f",
      x"b55709d621ee11838bea50bad9a8d4fecb314846b226bafadc3ff3bd4b4d19ea",
      x"db166fc1bc0dbe5208c8569b73cf5ce7b94993903e3b8d32707962034b2cd8a3",
      x"cb7ec88377c03a9dc8d08f0477e4e42d260165c75d908281b4e55331a5ff9d1c",
      x"c4e4953e426610aae6f81b22c2b57f748b78c3bad3d8e45bf52e2a83e81d828b",
      x"cc303eef848b3ab193fdf37b7da5a0901cf33733980c018dce9ee8bbf89de812",
      x"d6bae8c6ade428518af3264a6b8dfbd155abba4ab51d51c67930c0cd829ad28d",
      x"4144fb25065db15ade1b267f9281c30cc930daf6860a5b3ca5affe5e74e8433b",
      x"91e68bcaa8f2163a2f28ac3564c80cceb4a7f51044a5195593d1fe2d8f362a82",
      x"dc3611e93309ab23ce6d1d830da26ed0bfd3584629c3a0b6c1e29e6621c55fa7",
      x"5ddef800b5f029bee77626611d376738e177c9efc08d16641e6e433d3c4e65cd",
      x"fce772e6adaa0d51e6aa3df5f48132bb88dfdb01b8ca6af6e842d5300d6fabe2",
      x"f2f4a14421c03d7d1751da0845bf82e73f2c463789f0c65ee9d3094087a3131e",
      x"eeb8914e61bbd33b53278487666b5bceb7d58e0fe0015a11c694e96a481a5a5b",
      x"7e736412a6309c925a17bf859944466b4b663b10d1b9b1d71deea204e4c2efb1",
      x"baf9a83e400c886d87719433112be0f0c0fbaf3616f6040df72b997518e573c3",
      x"ff42f5377cbef99517f37f42f5ccee27076f4ae0bf8e1532004739c6a681562e",
      x"af02f3de6e3ac9ab68cd08aca62b6ed3f7916d2a2f0e846abe48ff779768e0fb",
      x"c526358501b494385e60ed8d08a040927195852bc7aeee35953a9011fe6e901c",
      x"24018354c4471d9291628382bddc5e1598f74d76eb6ef4c1e939cd0f835c2f97",
      x"64ad4d2585531c6b4f9eb0ffd4f6a01a5f957462f8803f59d48d41fa9613c45f",
      x"573f680904d0587f27cd742a9e6fb9bfad4c0d65790bc71aae5acc5c70988bce",
      x"a7b449adc5ca4f89b5ffd2f730a8df8dde2e7e256e7c74b9c5f53003f197f955",
      x"b2c5e29c8b345d23e9e88e9a9c11252e5d33acecd7e77713120d46a5a59f8c70",
      x"4665c516d039c271db8878e02b7d3bdbae44386761a833b006ae43172b618b90",
      x"b03e96bd05da4399d2841477983222793946b4ebe1380dc5193a50d02224b8fa",
      x"5b549b1f2420fb426c273b24377f516970ab0b229b0118def6a706c9f0c96053",
      x"e386dd81f0207faa4f7d867e94083b7d9974b3193bb3547880629c120d89299f",
      x"a0db730a39616f0320a68260e802f438fac3f5a68e445d81ff4a2f9cadb98d16",
      x"27d829641e9e99babc5d2a5b7e7db1125b72ff6ff882f519209207b3f3da2a6c",
      x"a2e4ff89daf3261450857319b0c9ab9a0c285d5a789291541d3b5bab5b91373c",
      x"e169529c9a91b8219311cd6fd3f7c8ed4b68d6488aac1b2d86170991386b15a8",
      x"4db60607b15073b754208692ed93c557ef8b1d7b76ca13e3e58126a0a90f3dd9",
      x"1064bcd1014b01847146fed28a71e4b80aeb8c55c2f4d7e7b53e353054040f51",
      x"8c71c2afa5bc63e9bd80ea3edae9e355529b9703094a0bafd4b1731208ddf22a",
      x"db3d3399958ce3dc9dcecdfaa69a0effb30bada61a4cd71fab3f224aaa3cc19b",
      x"1de90feace730b9d0167e562b95a6f50c1d5ee3126dac7109ae7d300a29796c2",
      x"48ec79e78f2a00d378569e7ae3a90d889d1652634b4c598510dd643481f6dd97",
      x"e4629a398d9cccb1e02f618d43b74d8e65cad473ac343b7a1640eab22a6ba10b",
      x"679c277f6260c373d14f6591d511776cf747720b2cf5c970d7dd3e49cb455165",
      x"80745d496e69d18055bc99840c8ed344b5896bf847eaafd409849974b97386d5",
      x"e84c0e3d5e6a81298f922452f4fe594b0a659f76da8d363821497e054986887b",
      x"b4c806b343cde9db76dec80710f3e7b31291fd455ba49a48e9dd74f97f1b35ef",
      x"38767e319b4f57459079b8f7a46ba5aff3b69e407adc7d03097137ec172046cb",
      x"e16ee502f40dbbf4a6399a052f5079a3e179437c3c3889d07fde5b9659eb296b",
      x"d79e1a4c5539b57c09b3aa872cc021c820981846185a473a0b74c70f2bce9bee",
      x"2eefa50ad5afe3e3c06c892200ffe7fe694a2db3bc2e740a98bc1bb26d903d9c",
      x"cb3889638088dc83740baf9003bd85823d7ee43bd0b34590fd5a7b480487e4c6",
      x"9fb49a49e4682c1a93a3c928c066c925a3414a4d6eb885d34ba9668bb7a588c4",
      x"35d74dc3d4bdb0f8571f518aab7ceb5ae5c53a9fee4acb8daac362f08ce81707",
      x"8705b107fda4e2ae29962de31b9590260b3f6ce20d5008139cc3b180846aacb3",
      x"3a4fd70a119da4c4716456c613ddb099e54161915ea5e2083f8982a04470bc7e",
      x"58e828d344dc752aac14c128aad546b194fd7248fb2a1e3488ad909e8616fc73",
      x"43ec125267148d616d2268944abf6a3122c5adbdec5cf0f52e86367bda37985e",
      x"f86671dcd5b515ef92915954d26c1bfb31433c268486648c302282885d66dc45",
      x"0c42c7fdf5e396f6fe2917d8668267d478442e5625991bf4be4411acb9664574",
      x"55b0fe76e75bc35a93fb44ba9d55143428893fbb2db9321920d97244c3a56b20",
      x"08d0f1df412fea0786c8c32826ce3d44099e0fb42bfcf5566af9ba5787594e09",
      x"9629feedeb89eca16a13ec8136c0be223298a5ec008a5edf543aa2b4c1521f75",
      x"f1b8f773dbf434537f4002359f35bb546bf9111fbadcc45b44d0a510af804eaa",
      x"e01bb93abb5b741c6327b819128188cb0005c97fb0288f73a22f2e62c48bc71a",
      x"aa56706e6a9ea09ec07575257ba9d6e65bf3c05cb4878fc4bd6c3b0c243f8882"
    ),
    (
      x"d4b9bc48fc0888eec5f8332a54ccfad9ad3e8e3cf7735db63730b47d8915b173",
      x"0a2c4422c05df99ea392c033d721d302693e5a3bc6894867fc4c8360bb9e9234",
      x"ff1af312b0fd461419d1187b583b2c0bd226fba2b47a72307bf52fa39cf0f37a",
      x"7c2c2b5207bdb39cd15324ae91f5aa77beb726ec55a198c8291c0be23db0d291",
      x"e284babd22bbf1b9c620be54235d7f62fbfbcef1268efa176b7b4d6725f8fa3f",
      x"02eee0c6b254d2bcecda2cf9711ad27c7af21b72df9dc1c572c3d18b7cb94b3f",
      x"3a0b40345e5e365d265e4f6d52ae1c17068517722a7a12733072d3a49a6615de",
      x"a3e55dff96a2b5dbe2e8bfc4c9cfd84abf0cd1304aee59509b35591599749816",
      x"8d1b7fbbf9e8a58c58fe3ccaa5df28af4a91569c3826d81b90404fd93d18e176",
      x"ac97db21b319227f6a577895330588f123a361f2dd5150d935cd6f8b8cac15ce",
      x"c471db2162c845abb0d23c32cb598b0b7bf1daea211f0ee7fa65f330e275b819",
      x"e2beed268273f3c4b4848906ab8d0d3a36b1fd071f3f3515924db7514b163428",
      x"c6894d113adfdf798061f52085f1d0206d82b5bc37ca34cbfa7e7a29daf95733",
      x"09e82ad3a5cf93c38cd1cbc194f6e4d5e7d8c9cfbf11f4ffd5eef52b38283971",
      x"ce72eaf5bcd0b4ff36be6389cb176d82bd0608335bfcd0174c7d1e7547abf4eb",
      x"0f054f4377e4314f15a51463c167c8b9de61280011b8d3398711f2457489e909",
      x"51835e56bab7fbd85663f196acd510c58b483ce25f75eb5092c7681a1aac7f84",
      x"b3a7069cbaf95afd4bcfb35c0de8a4ad1a09ea3fc2ce61a6dd3c2aec731904b2",
      x"3bdcedab0a749df1d3754533c4cd0b4dba6feefc06263c2f418c8ddea029b74a",
      x"ccfc7fcc42eb3926f93a6d1bd8fec95b7c69e2d7f1448119cf17008f9e34e10f",
      x"a21b3d4a3d6abe03674b60cc35fdaa8fdd43b7724bba25057d54da5d9f8ee4b8",
      x"37516822b15895f93f7a4a726de4a6c5b30a2949df1d921732ff8b274566f04c",
      x"b6f8cacbba9f8c6e36f9d27d41a3d217e06a4ec54fcbd32ea5a90b2b83cfb40a",
      x"7e180db46396f39d94162ad7dd921b72952b4a2312ba2ffa8accdc123875aa45",
      x"73607f73069c9cb584b0bedcabe53973f8410b20e554066366899a6e353cacc9",
      x"eb6c8fe235e6a6c9d58d9872d67d44935ac71a800607bfbece54756d276b6776",
      x"fdc46735f54f423848219588e1662893e8e7281514227777ae4c982ef92930c2",
      x"7979fc070348e22f5e470f66ce264a8ab401f091a8c060a67fa210c48e3c8154",
      x"aeb31109e436bea8f2d4bd4823cf35ed2fd72d7afb3d2703eeb20bb043b3af23",
      x"595164ab460c705f059cad9101a66124165ca410180d90eec1cc6f35e1ace1d0",
      x"c110a8835c63875d81b8876dee5c0aacba4e085a99b027c151c97bfc25c423aa",
      x"f7af622ec1cbb1edb0b875250b358b94c6edd40a3c068222c9f6c7dbc2fca84f",
      x"a0983fc1dc9a16e8fd8f4572366bb6f692afe00e161047ccf26b7c856be57fd5",
      x"80c5cdcc398ef876cb96f6db2de674e23d0253e93bb880e8759a7dba05f98c71",
      x"5cea382f5a8593a2ba3d920525369ef40c778bd798d1be967064e532d7d68899",
      x"f0c2abb52b17e29555932aed5ccf270d563652b1f15584f51fb623d5110cda48",
      x"ed46b11dae5a97b567fd1116ba4b9cd67a2e1ad7482c3f25016234e25a3a6da4",
      x"7d6d7afba95188536b121989b29eb7facbcae4ae9298717a9140cc881dc64997",
      x"21436a9f25ee9dce1d7756ced548f4e7000f2802662bfb6c236666e6630eb9d8",
      x"90f49b029c740809d1d6484c00eb41e0e81bcebfb4df5820c5797ff44e88ce22",
      x"abd4d3888f997d033d4d64562498eb580be976bd566dec77810cd36e12f0bcc5",
      x"b9045dd22cf93805592b2c72813aee835148425ea5c35cd2c27ed1862c0211b3",
      x"afbe4156951a4908484994a35f5fcab2cf8ee7f454e6c1fe93a0566a15a0e07c",
      x"8a122e10a12ff472bf068067e8eeea16effa5d5ee8ecf8e16389db2fbf9a965c",
      x"dca7abca0094456ba8b7244268b4a799d4e45059a6837e2f47e8f086f345863e",
      x"ce9ea6ba981a81a1fcdb8d60d6efee2b822f936da1971865db7d3948840955f9",
      x"b4e9d338aca4c9d17637c0dc50da8e554d0c1b74750c99316522fb7dcd6ec5fd",
      x"c53e25e2cc9b1f815e24f04195d7128c62d0f9b129007fa8165c117ea4771156",
      x"f90601f34a721a7acffb8ae0e0d3d97d5c66eb1999271956e1129935ba93a9a3",
      x"cedeb5a36ba46dc9fe375c945c5d92e42fbbafa77ecc3ea15a23548064176079",
      x"7ba5e47b3be1279f753909c72d3d922faeb7db070123f4fcf3db98043bf7bf39",
      x"3771d98e56f2869593a22410dd993ea1a63e76a0962ca609c59da7b2538b9034",
      x"d26c0f9d2cc308097e67ec71fb163e1d94102a98eec97470880081fd43c9264f",
      x"db0ea0af642d16e6cfee0ed445b9b79f79a9d7f902e0d97c29c3a2f8cce75499",
      x"393e13ee1d58d900f8ff3d19000a1f2d99abf58791e97e66285cdc5819f9bac7",
      x"af4ee43841712576166d2c85abe14fdc9631e8bfe96a9828b7ec291e37b22e51",
      x"476ab009dbb8fc2cffba93d3ab5febd09b8654af4c92e4a6907b8c38c9bf22cf",
      x"153ddafbcaa40ed8b44f6967f5984415f8d7ed53caf9b497de4ed6871b524ef1",
      x"b00ec99b3dcab4dde16fefa7734cb103b6918c1e84896ce3241544024d049ec6",
      x"c1e7b63922ba578743bd676e54da7a798f65947d43574709da9a60ed016990a3",
      x"601501dd4d39728e40c23cf9ca6ea69cbfe401eb87f0375654a75a04149430f1",
      x"53bb016dd8fd7aa73d49910d4a7022dd063fd7c4967e75cb4ab1327d66fcb71b",
      x"08ba60ab1ce7acc5e7a6c535305ea26d7eb31be3d70e91e353c7cf97725aecf4",
      x"21ff6d1874d324eff3fddc97e4fddfd494db2d9dca55e31af5431b0a39be003b",
      x"640352e0af1b7873301ca3bf0a6d8341d98631e58b34aa14e4d81a3e5a87adfa",
      x"ea2c836c6cee762dff75a4ca251484079aaf434726efef69d6c05d1ecaa08884",
      x"724a9dec03eaf4469a00bf7188ae14f793392559e959bc6eb1b61ff3856dad5b",
      x"ce6fcd69b38677c477dcacf6526e4ca60c2704ef757cb8cc9ba8bb723b0b6631",
      x"18742e39f444d50adb4e0d08faa1b16808e7559e5b8fec9ce7bc451458c61d06",
      x"54fff0e18fd124e231022e10fa9137140bf502ccac94f9030355cd2c6b031c05",
      x"979d0916211429c7bc1911fecbed50d6cf1b84e702f498e1e87ae0e92020e267",
      x"ae5caa9d26e7300f4e38708e0f91f831ee87e2fc4ba2dacbbd8c7cc2e4b33532",
      x"b8efed172af27eade00471a27590874a5b4db424c96f14db6c5a7e7cdc469464",
      x"14a8371b2fb70947add0d9efc8dabe69c90f058ae186ca31522b2236c7cb0e5b",
      x"48756f2ae4aca62956ed6c5e5a92f9980328a666fa1364e71110a540364572d5",
      x"c8d377d1aa7f2d0fca0714338ca1a2e72767d0b0cde8f55d852fc5850865e54b",
      x"3d603c1335600ebe918f39bbc3afb2e63cb0a2abc168b7d5c88ab2e74b8b97da",
      x"cb643dedc1d34a1ae02388c75b9354d2bd7029688eb8961cb93528beb9e4cf5d",
      x"ff83dda36cc3d4c6f2f70285ed5df9def7df0962d8902a91f1db70c8bff08558",
      x"0c0626af54333fb12ff7404fc180485e131c3c82505c10f61980a40d60f94562",
      x"0de145d6768a5d27bb81ac38d271bb7e80c180c6e56334200bb0c77513d7f0fd",
      x"ed249a567068a1448a76cb4118251727a02e60252656613fc9ea42bbeaa4cafa",
      x"c4afbabacfdcf7b616e07ac129f9e70bc357bc3c20fe8a4cdc7fdc4f65d0dc78",
      x"d237d7c0da4cd4c5452553808c6c34ff7e69d1512bb6211635a927ab672d61c2",
      x"ff5cb1db8532200e492a80905bda6903b45386cc98a74bba24effba154e4fb6d",
      x"cf3f05b7085f009b4675d163f83f8a98d2c51afba36cf43489eab3f1bd56305e",
      x"e8b242e89260b255f5da38eb06c5d76bb353dd65dab5c1d20e4afd0fe36e19fe",
      x"42126a6abe2125a13d8580392bd6eaff56de01fe109420fcb35836dcc08dfd61",
      x"67a6f0852e252036ee38112ccc773006d2b7fce6724af083af45b20fa96381f7",
      x"4ea42e44dc990a70a6949f39306221cd9cfc80fcb296d93b6393db1807daf0c0",
      x"00ab57e860edff9ec9f747d5bec5c9cdb96b86cc5a1c3a7532a1ef528eab222e",
      x"45498cadf9525ccb056ad61bee32b8e00f97cca5cb040131b87656676c9319c9",
      x"aea9cbf1559232a7aeb2ac53ec9407860dad3b12274c085cc11218d5cceea525",
      x"9d6824e5d20db6b7eba54842679377f7f3477cf40c1ed51441634d5b8c16f509",
      x"e49a43fad0c8f5bfd59e39af7b54be897a70ac4983cdd0176a5d6bfd7d010805",
      x"c7273eeb2ff2c082ad35eb11dc2ff3b79cf6e56d06ba79df490a84b65bc8365e",
      x"23ed10c628e2eaa845998248daad8e28a13e940ec56e3ede74a2861db25c80d5",
      x"9ea868168bee01141e4c5222fabe5119093ed41a0e9491327dc935e22f924eb9",
      x"3f0ec4e2e8b5bb5bdd6befcb87fd4efeed431ae91d172caf1874626b185ccf69",
      x"93c3ed1ec607ef3c902b515817ac6d06f7030b6b7b7116eba9c4350780ce9ab7",
      x"43c502e538dfac60d86005eafcfb2382ab325192de5cae10848c61a9e2ac6802",
      x"b0ac0d650eabbfbb64b402e7a56859438777c5b8dfa35a588e713c8598f1330f",
      x"8f33d51e2412b3c6ee3ce1807ece923093d78f83b2809c37ca23186495f0ddb9",
      x"f036e3ebe71b9f2b1e6b03c26c76454a4e04340d440767c5556c1e04377a05e9",
      x"a34979e39c6b768306a2921c8188edfe4e0c3f469bb753870cd2c933d3a545fb",
      x"8e6a5d77c20c3e137782cc07da6aab10984a491771765899e0beabd2f4bc24ff",
      x"dece568b39e62a1d31e5ec834a9417566979066a2dc953221cf13ae63c1c881b",
      x"7403fa06b4abbb8216534e216f306caac695bdb5153e6264f971b20bc86c940c",
      x"3f51b47c0136b7efd51c1e2b425cfacef22c79a3c9ae6e646845b250725d19e9",
      x"1401dc690cb5c7961165eff9af2acd7fd5e1c7b05c32150d8392a8f473fb232f",
      x"3bed121f4090f01cd5e0858569ef7d0b5181fc934a0110e7a3590959ef91482d",
      x"990d3be6e3ad0d43dab22eec6a1ca369967b0f45121c4b423deb9ee7f7e72acd",
      x"737f6d46da723bf249ed1745c25ab1fa28f702b9b4d2fdac9a42e1dccaf205aa",
      x"db8438dae37939ada35a16e50279fc013b9691b0be27539bdfed84dd402e58ea",
      x"f367090db9e60ac8d01485da2cb910303458dd3d36715fddbc56b95ba0e1e483",
      x"06a91cd77b242c3f3c12a1d3a9e7e5a4132804df43e2e841b000ebdac23ba859",
      x"af33a2bb7a17875395958dc5109f82b43353b1417d592acfdb271115efb80f30",
      x"c6f382aa4435482e0b0bedf4c32e2823337e310ca1d38d1d629a999dc2ce15c3",
      x"0adbad8aca389ec562aa4c94264204caff201c4a604c9901580866cb98f3673f",
      x"da86c4df8e386f5f47ea3d1c0c451d8ba6585451d8e891a2b69bd26e208e7cd0",
      x"4bbd9eae9d149b45a2273e4e35ca5a5616199339b18204e7bd1bd3f3a306f96f",
      x"7453b30427c6b3a0148ebf55e7be03c6b53d04a2d6b8dc6608bbf0f094bd5336",
      x"ba24f18c019a2fa719c0c9f66baa6b0860f5d060aec13adca7850036b2cb8e18",
      x"d201389664d269c0b8e5f6b153de91dcef94e22d4090086c10631e001a5c374b",
      x"bd3d149cf578dcdeaf091798e4d944ba118e03ade3393e25222cb4f5f2ee4912",
      x"73e3a056f630ee74c82c6c1b0a0ead486ff7bd3d9e98afaf954ec05540634d03",
      x"89594ca5a3be567484f5eb53d69abe0a16fb13a78f5027f36b059eb56fd7340f",
      x"9e546a7098da56863fd9f76678264f08f1bef019f993ff4f30b3d4db467949d1",
      x"a90e2b5b9f86918b0f2e00b02a07ffa135027b310107407c206f25dc5e82e766",
      x"a4104e81fbb4174fc9b82bbd79b93e40e0f89970419f5616e9439c43761c6bdc",
      x"24aab139ea642828801ced1bfa44f3f9c5277d02432a5bb4d5b22b3bebf39a28",
      x"30b2b64d051182e99aba688ae674c20f8cc44dcdca2bd2238e4c220ba1ded858",
      x"cd90739aca859a27e6fa12e617a9e4a162a3b15b355aeb48de8fc94b459ba767",
      x"36059fffb1a8c0426330444fcdd7b35748d4d93b41e208bbcc25bb0981662660",
      x"c787e99b4cea2746b5a859e9261a2850124dc64e622dc51d8c2710522c7553ba",
      x"2eb3750a9f804d138674abb3757b63f08ce0e4e61f3599344f2a9a3ec79967dd",
      x"db1ca1d8b2155ff112f7e8398f70b15e2adadb48538b5e897f270b1c06e4ba81",
      x"f10075948f1c3ecb46a05f7391b031ae3d3c356c1a4bdb4d961bcbdfda259876",
      x"f81788f1fe8403f290e10a1b84f580b15ded43e1b3a2c8bb8de9df863e276f1b",
      x"84eb677f199d8dcda7132f7e780f0f99e83bf8c45be9c5e387989eb7f6b3f225",
      x"c88fc57dcd9792d1074088039b707081798b259b4a3626b9fc3f9c4cd41d234e",
      x"de57d01760cadde8d08eeef2a52130d552f4c2dfe80ed7dc9fb55db295933b74",
      x"43e73ebd6906a0bebceea619b9dbcb998679f1e7c3e41ee0f5f0cb6fb39b43bc",
      x"fdbc363b9066848d77ab850e9cb0db4aff2cbe69c532a5a4cfc3a1511239be7b",
      x"4f9d14e0cd2bbe2c016c9b62b5512eece30a5bcee67c7bf2e599f7be6b082bc7",
      x"a210c84053a85d62a2590ac84d85438a4ad75a543ea7b6f1961150098c5a7a3b",
      x"b4229a43de2a3a18fbf9772891e98a3ccbb1161ba0e86839a4b9fae153b57565",
      x"4d48b7c63861722ab9945e02c474824deee906358731458b339beea25756170c",
      x"ca9ffab49c838c638e1878d613620a0065e6c4e68d270e8b47d4eea9b8d435fb",
      x"88ab5330da19b097725569e84e7ed1febb181fc1fbbb723bd78c6d314974c48d",
      x"b2f49c166c4bb4fe80f6b5f0af29daf5ce2936099baa008b1bca426567000f5d",
      x"624c7f9690750417e0dba2a0d213daf22feef8f6d7d6f8551e15e8a17704db78",
      x"723c426c04f89e10dd15094f1196f0b9552c8d065c3f063e16e677fcffc1a1a8",
      x"ece1e8abcd47c472a24b4da2e025d87ce852092ac35edd9d2f6a56e3d6f24f8a",
      x"6ceeb11e19933f0998ab76a57cf6b527113a06317e1009253f1dfa46f35e0cbf",
      x"387c85653e8fd8b3be1e862c5251135a077388b70dc4e80f20ca692133b5f14a",
      x"574b34a2e3b87fb7f879df014aad9916adfaa3e7eb25e7a2c044b59964c6c970",
      x"325bc43f923154f3712d624a0dd7c67ff72fdd5be7e2a9f76ba91f3e58625ea8",
      x"54567ee0586ed23f9e4b605caebaa2d31b0c13526989d03e6d474f37e815a364",
      x"49cb675de9ac77a3dfce304ce5bf98a6ec49260ba39b72b6e895320c3cb8b4fe",
      x"f2cb8aa1968d3d50e96a7c69d538db7554da6a91f2f793e0c054a7c8f3c00f43",
      x"8d092c06b3e5337c3881b1792d158c6f053baa24057521081cde51fd40abc970",
      x"5f624fcc7cca401fa535787d8bb7aacc6856584ba3aa1e2fc0caed5de41826fe",
      x"b416059b474e12e412d5729475724ea11587582a93d82f938af570a8de3de4b9",
      x"0cfae5a74627eefcb6d1779ecfdb51372c6b028519244ff6f94e25ae695d60e2",
      x"3262fa8cca52f0c884255dfae3e81d5559d1a1e66858945ce3af0e4674692ae2",
      x"5162f297e0fb2d8a826791ba1f9ea23d4e65a55a77c67c0f7f8c46cda083f3ed",
      x"19b3fc5bbedbb6130fb4249ee7dab2f097c98a27fb4916a369966c58c9836272",
      x"6b2ee6387a5537b199cf29b8f5ca4066ff5066487f7d28388c2f3286fafe55fb",
      x"b71073c12d3ccd308a0eb06403aa5b1446dfa6966185b8369b5894d72834fef5",
      x"c8667b59a9f4fdf3e552037b9dcb9e1f597985fc8c470d412ecfdc35c79dd374",
      x"dea83563c82162eb25bb06bfd13846a6b4d4f1b1a7137bfacf726ba8ef4d6fbd",
      x"a50805800b209cd49213da539ac50c355ce280428a5c28654773d090a8f0c491",
      x"018da79e8554c8c77875bbfa4461bc072d1bd0cfd39cb95ee5e906021ce6a784",
      x"bc4a817cfa651c70a090e260a518699ff6ff5e066b2e2f9c92a4f783c41a9abe",
      x"602924bb307f41148a6f1b26d391fd9a36a609eaaaa6a67563d57413bf7ce833",
      x"009716ee8695811b7d7b3cd2815894b3b8e1fb280e4efd82f092d19473079f81",
      x"e1648e7c33188ce61bd6caf50aa67762bf185c622a6ee5a05cf40b8a3845d1ab",
      x"88b18b2d56e90d383da980c31c00748a0c7284b3dc90179b013d5e4ccf3dfa6f",
      x"15494429668ead8f902700664bca2469fe4d4469692e0f861e95a3982ffcdee5",
      x"6e34aa49687d09e066d7758f3b9cd0eda5e9305cf037b4fcd988c7262d3a12d6",
      x"b6ec765652b447396a4b77d05e0e62e0050bd166453b90a0e8d2a4fb450f3bd0",
      x"07513c580d1662b7322737d717ebda2e67f2b0f5bea7d81a45b85730234dc659",
      x"37093d1e68c560fa49e0b0a12716c4aa2eef5ed6a8fda87846c2a51e2f0c2df6",
      x"62939f04bed9f7501376157d5238bf5cb320fc1dd5a30a26c3e251156adab874",
      x"1a33d5c4eb1bdd66a4ab0635403583b36e76bd0c89967e0091db99812e858cb6",
      x"6236cf5044e59ce74fb53aa403b1a7898c96d7085e79810bab58e4601ebe433d",
      x"d7296913a51b999dcfe6cdfdc014df658a7abb7be12b035032fc112275555dda",
      x"c397a95999e9fee838bca0c11241a9772321544c086c739d03939fefa85073a5",
      x"e1f9781e74cc81563b100c5c3e11a188fe623a90f187102e3621dada14fdfef7",
      x"14f4415223adea4edf882ce35e110cec02ce61f8a72ea3b27d8665d1f0d3a9e7",
      x"38746a1f87db291d298a79d671a2789cf3ecfb0f96489993fbfb3caa7e5c85a6",
      x"ee6952cf621a4de1d372b2d68bcec6fae0f15db5c41bb8866fa7de6503935172",
      x"41b2ddbdd2ac4a3d204fa094ddc8722f3700262ccfa4dfa0f8cca6a22c39f9a5",
      x"ba1a4c2cba1068928f285fd6b75bcba711ac573f533ddd3bb468ad6d388ca577",
      x"c7454363639bd03da29914f18b0033b9735cb1d4d5e268a7b1d6f027e742a207",
      x"b6c7a664cef32eb8753259b7de6435c2abf5925390733bd4d830eb4f6dd2fa60",
      x"0419c90c6689d41f9f8a1823215370cc5af64f1f7a168c1517ca6ccb4518a643",
      x"0c4caea459bb930d4969b35bef1b378dcf9035881372be46dba7515b2f9f6630",
      x"fb91484c55b4c8c58edf152c4005ef7125c3021e6f19fe9edd6a1dd231d93983",
      x"4c02cfdfa319b88f9d1a6ff65f0f62b933372b38a0530cdd9d10ad39df2e8eaa",
      x"4ad65f015c26cb69f0994b3fcbd25c24e415cf2e1a6ef8d4b940aa8e7eb5a80a",
      x"77d5d79b9ed9d88aa201d0620b173be7ecc9a210f68c8f3bcf1f0d63275b7fee",
      x"41d7d18e5301a456d97b0f6951554ab03e37437aef6e8ce4afeb4b0e6d69260f",
      x"f02128d59d288926a66357d9c9ac053a483ebc83af179b76047fb6b9b66fb4e7",
      x"b887b863c9f43d0d523231d26a33ededbf62214bac71dcb67787b07bd472f797",
      x"de460ef923cedf51f41181a855dc64167b5213d6dbdab1e523952d5d8e5a5ab9",
      x"47a7482492fbdc24fe1ec382550d4ac509883c03373f86307f57e19e70e05325",
      x"98f4ab28e1b99a48ba4f95f43f5a38baf6825e646dff2d173df02651514a2709",
      x"7cb93e941fb0e3f343086ddb274a2c3ea50ba9ecab20e8f9abe5289ae65ab146",
      x"2da916ad096dcf5ace3837daeb8d0aa0ba4c1b49f360cfa108d06eaed91cc32a",
      x"d8faec8ca106a7150cc51c9024cb56709c5ff13d9c1739653dd3e49fb2ee71c1",
      x"452a854bc7270927854a5afb37f84db38108649cefab9dd678ad2a2f00a2ea70",
      x"03d35ff0e30ba43414f8216896c168521fca808892f86eab225339e5d1c8213f",
      x"4a043775da8baf5714c77da87666773160804f9544bde78f811228d1d432d121",
      x"4871d9877e4daac5e151580704b2191d8af4b313f8fdd3e4d1e0f55e0d52a1fd",
      x"f5f10df53c2b649ec6039ece5e14b57ff055970e2454905c7a28c30934e69ef2",
      x"7ba53f810b0eeba013f067c32085a550d9e4cdb2b0ec422330411e129b00bab5",
      x"3deb5327b1f4c6f6db3b23973a93eb458560f1c4a8838888840bd5896aaf0ed2",
      x"717fced2e4750bf4fd31a5941ceba560bf1de5a39a4c9ad0c6acce171c9fe257",
      x"3d03597f2bf17d4960f4b014a859c90dab9ba8cbbf244fa936e68d3a79465448",
      x"30faeeb72f94081b1e12d53311d558c1a6389b39b93b3aca0da973b8b82348e9",
      x"fd42dd70569deb5f6eb2cd295d68724eefb0fd5c6235b5e0bda3b1ff12a5edb6",
      x"4493f8c9fc884264f7ab2648b1056f8543af632de210c0e4b5e4b7505eedf726",
      x"c803bbf20d27b67f4e3de1075c1e82e442927e6b439c17cb3dfe3170d822e1e4",
      x"38616961229484353879c3e4bb9f5433288520c184b1d238cdd9dcb3d57ffcde",
      x"20080febf874f2d5a0fd4bfd80940d29249f6bdfc0411ebf25bfd0816b993b61",
      x"866e9b0a9776db2388f022f97ad670f02a1979da11040a4a30c0f628c0d81217",
      x"648cd3323902976ba4dc4dd76d9c1da768af1d37613577d3fcfc6a7499922cb8",
      x"59187c8976a637e5476ec77bdd773ad055b79aed92a5140516fb9b43765e76cd",
      x"46d9e8903f9936511f28ac3f02a085669708482cf6cab83fd33bb754f68abea9",
      x"ac20585b729caaa54f21450cd294a1ff454f42f312943eaf64d6b2ec8222a479",
      x"99481112405a447eb68f08af3a6e5bb38d688922018dcb2ada2d30ad2c7c92cc",
      x"d2d61e2e548e0361ebf799d973ffad29cbf59c23ffeaa86d94942eae4a516c70",
      x"dc8328a80e93e53c9e0004b6b4343c45460d072bd178cfa970a7175786015090",
      x"4233e9c09ce7038b3cdb723133ec5ad64808ad656691c6d79a49c8b95fdfefde",
      x"53ec2c2c90218b9911b4f927c6a2deae38558b27735313dca4b69c20da723ec8",
      x"276907347eef94f25eaa4741683895aefd30e71a6d5c5bb847b184b0cdd544d8",
      x"cf40cfef5985c7c60f8f78005e51e59c692f8bc1e9b8fdc93d029b739400412d",
      x"684da17c290d108b2d4b0bbff785c47e82b26b2ba96f45ca2e99f3d6ad1bf8cd",
      x"c0fcfdb4051fbe4a2608083a2a8aa4a798ca8821626996287df70bfe2760cc9a",
      x"43f1a783787565b0a8176f633ae2018efdc9058a8abcbb0ac968a4bf085fabf2",
      x"dcd8580335a78cbecdc16f4e14f3b6ac913eac1e5df266ee089fea256bb9d0b9",
      x"1dd359133941ff6d93b7f2d6344dd106b5038d4c2b08f59e96ab52ee7554d67d",
      x"ff80815d5ee613b39bf80dde44b241a1de858d2025edb6f52a06814bcce4e044",
      x"27d7c48e88087d554f4a63a263b67a62c20df15b94c4dd67028289fa5c549a27",
      x"ccbbbba546098a19cc690256ef1d5a5aa6fdb407dcb0dbe5210e93bdad2701c1",
      x"e359e692fb58b80b52b8893f89b66ec6dcca112c67ca77255bd1f125c0b08eaf",
      x"e231e47ecf8a65eb2f5d5839c98f8b4ae7cdff4dd87da867be84122e64a6ef08",
      x"98858ac8b2b1e4477b21a3202dfdcdb4501b371f8856a63bb81b6384019d974c",
      x"06db95522c16fe4ffa4873f663ed9d25bdebe46956e2206c4ccd4798cbe8ebec",
      x"44ed6f93f8497e66239685ae99e4759724847bf6f60398b631ff2c1103c43135",
      x"196a87d51ffe53041b2a601d0de3c4574abadc253113b6552a10a50735f379bc",
      x"71f442e9ac26589850e92d40f189fca2fb286c386f53a56687b9b680190698cd",
      x"32c13e5ac412bc407f68144aae59955989b1075769089bfc47f08d848d7e2d44",
      x"18e848d4886902f50ffc47bc7c2554173c26522cb0a3445dcfaa37b8a1465a4d"
    ),
    (
      x"00e5c3e685c3f6a8ca201cc72d539acec8cc07ef28c72ecf5d901766cdc550a8",
      x"3bad4fcc772adf65dbdb88b4c7e98867d31db754bf43c171731fed8aee5adf05",
      x"c515cf64ba9fde8db31d149b6d73a7b3b777ff33de68e7bc6088c1afabd241eb",
      x"d4d140782dd7c1e7e57b0f01c053f957ddd1a2939897d255a6b4607802616f13",
      x"1ffe3e82e4fe9467d8d6f8a3b97c5bd5c0da81d3307f2d19527a3307339c321a",
      x"ad3d04fc763f4c4864421db0375038a93dd58d1e0b53a12a6947240918040b25",
      x"0d8a5ddc1244135493464dcec393966c653fa2e9de0ff91da4355bde60e956d7",
      x"4474c494bedab65add09b4e8d8605d4b60ee8278e6962e79d206a0d51338f707",
      x"254ed72be46a43bd855df74a8a7faee5e4c79f7136e98485cf1a7df9ac7feafa",
      x"2f619e3a02b26199327ea3e60cd785ef1bbc6967e596c779620b05a2b181b6b5",
      x"2adcc8c5ae632fdc86be6994499ee9fc2fd412d82a02b1b9f103c8ade0307f5d",
      x"5edebfc0b26798e1f0f85239c8de2f3ffd39bbea9a4e166ca016fa27053ff7a8",
      x"3d4fada9377bef80195e04fe544836cd063afd99b8a43c2f32870a342768f952",
      x"d7329beeb64ac413ed4358e368f170d7541301413a11d15193f44f33f9b7e455",
      x"9846b75825f1c912fa36b845761f7311f404f41056e8a7890577c32ced863e83",
      x"6a462eeb6f51ebff947d540c407a95ca0b9ab1901d442d00c579db6fcafdb3d8",
      x"da7ebb4e58f56f19df3f061411871420ee04aeaca2074133ab33ad4311d96215",
      x"ae4364b9a5cc2cd9977b867d8e5b55b8aba8e5c1184a4e9faecfc34dd7b290c4",
      x"067ae8c8e2ed5738cb73e618a53cfe50e561854ec160e75a88fe269529f80048",
      x"3132b7765387786f366539480256197bdd5517a83de9328b4656baad4aacd699",
      x"8c9051c80a4478b8e32b4d42aa032324c6c1021aae2f55d634c9b2dad15f179f",
      x"190b27cecd31c9574188b019bae9e8adcda13eaa118279b3933a89fd718c847f",
      x"edb799e435c793313e5d357beed0ee251646e3a48819ce4d84eb863465245daf",
      x"2deff255ed12565307589f06bf8955d3e5fd9fa7d8c3d7cb1843cef4ac1dda0a",
      x"1a053a10cc9ab1197463499b3229be12db4b5b5e0f759435ad509398b1b1400e",
      x"5bb118621dd14488138336bd3b0f4ceed6924594ea1127a273a71278da503277",
      x"6249a0bf8d92b3ff867f08122461e3953829136f19580bfd9e6abb01a911ce1a",
      x"24ff19e842f5c7f70aafa7dceca2e13c987760dd21e22249b81b3e97c6645237",
      x"8a1144d2b0e86c88925e133c06dc1da3f1e0f2ad3e9ac6138b5aecbdde0fccb3",
      x"f444be7966b10637ad8d3277d48133d01cb0e6f8f6bbcf564b25a72fee7f906e",
      x"1138db5dc62118ee204d03eadb7244d1a85042bf50aaff331e2d29c90c60e4d6",
      x"88ab6a21755572d81cb2c48bf4c3735dc04e67ff3c28237a250e210bfaa2621b",
      x"a1c5eea1575deb14807e19d80c9f0061ac64f1ba236d8b15062ab8fe2b276d92",
      x"2dd8a74055910292cece5c4a7cf0a7ef337569a7dc327e0aa29d2e76f70c98ae",
      x"ba0ba0c0f82f60f456352616ae2aeab013ba78059bc72dae6ccc1c5dbdfddadb",
      x"886075940f45d6dcc0519a5dc404cd199f2f4c2fc72ca82bf7eb20601e867148",
      x"67e2fb971b31f65424c48efff872c363b663d80e3678519cab5c1d5edd3d6f8c",
      x"4d9f21c82052da5053dffc4f1f2155f510d873da87abe79642f28c8dc6726c90",
      x"c412d73b6201b7a5103de2fc660aa0395dddceb70369690edba97b2b7e0b2ff6",
      x"04194024f9af051001876ef3f6f939a3b2d9e8b5c283dc5039e3f3d251cde0b3",
      x"f8ba529594db76f609c046b2a15f6178d7ccdce42393ea6c804dd3fffd272d2d",
      x"38fb4ca3f631ce555042637dc6099504c3713fe436f91e6ac20b496eae0f9e8a",
      x"eb09832981b48cadb86289ba5513b40077283638ef28952c418af431fe4335d0",
      x"da9c325a32a1edfbe454c136227ac53c539e428c12ef66755deedad767f91979",
      x"e1cbd796cb0195cc947bc7d7449c4f29cf0c81b4acd325ff8aed0bef0fc1fafa",
      x"b5c3cbcd28348d4484326b46194b47dc00bed00b8f012c6c02d0190d92a19d02",
      x"fcd701caff57bf5371d22aa229299c0f1b99aa50fbd7f50247038cb728c56e3d",
      x"9d0ff103c535b4c06ad57a1fe91f03d90e6f342f5bf1b25f31247a865381d27b",
      x"b58fb389c444635d7ba163d02526deb22b6cda7c53f76f5e40876591677712a0",
      x"64ae186991bfef514750f92ebad6dd4f27638a26d034b3cdcfc3a942fd5d40bf",
      x"badfd26ebc912bda9b747b84eebaa5026f1a95cfa75f89c979c4b8f10b19c9d9",
      x"70c8fc368b4b79f273a99b49f55f0045d922b31849445665cd44a43d196aa6ae",
      x"74a6e566ed7e116881c192099f618b5aaa202ca630f0e5c6e27d51b5961fc1fe",
      x"9bc822290de4105141b252bdf68c6d2f3eef26849b5fbcf1676ca7f302a2bb81",
      x"feca68c603a1f98c5785e0063de34cf03b7a039e26f011abd7151f5cae1075bb",
      x"8b4a20c3ea86b098c9d4064b40d5f6d0511af66bd3007c41d6e5cd91282009ed",
      x"cd96bcf17d967ccc4fe4492f6079b66ab64d3267faefe46a2537b69bd930b53a",
      x"f0251a5c1b86a7cd0b61b8fbcd8af790398d755752ea370aa23dd1a29a699b6e",
      x"58645f94f540ab585dd858d372c4177e4c2a2aaa965b64661f1d3f1002b63889",
      x"45626764809c1d85a50e3a4ac10e65536c84ba303055b11b7e27910bd1918abc",
      x"155271b38fc9ca156fa9eede1ba7088aa4b8c1d3bf14dc2dbbb33ed5f45b1275",
      x"65d236c43f1b39a605f1eb1db81dd42ca70f1f3eb45ec8358f7a424d6138f682",
      x"495bb7849c03663e1b0814b2ea7b5b88000bcb3b3a5bab4ffc75536decd288af",
      x"3fd1380aaf02ec909849b74bc38c6a3a98ceacd797befbe37097153d56ec05ea",
      x"dfa7b432cf6001446d9ea0b954e71be28fc053c55fd2b223768b81796214d472",
      x"e60532ff644b515c9585fcb57ece59386247366a116f2e63c04497ce8a5b81aa",
      x"33ead2aa68d1dd28d4bd2c12118c1867ad439b78e7b9d321216cd5db2ab24884",
      x"6f660e88182f1ba1fac22ecfbb72f744ed749beb1f09bb8974884e279a823a7a",
      x"39409c2ac05c914bc53418a40dd73834fd453e822d261e235fb7179de31e52c2",
      x"9ec62d7ba5efe48b2efcef3a208dfd14c7601a4bd90058a76857d718d03e1587",
      x"23d86cea9422fdcf2225bad8680622876ef9bfd55bdaba2a8b752ea56abe4884",
      x"d915e93135a166186950fe1f53b30a91c1327055e39b83d15aa7097839a32d67",
      x"bfd08425a7103a9d3c297378e17e67b4f98bca32e25f238649b9771491c9a39f",
      x"9d768f23afdbb763ddb0e03e2cfd1c54546d3331555ae3539dff41869e909c17",
      x"3eddc4fe8c0c32c649db93da5ab9bd8cca691757f01fdfef73eac263b7c28f55",
      x"6ac06211f2d670967acb0146bed8643e438bcf02460a32aa70659a539132f6b0",
      x"4b1e15987e39fe381e5f7833fe187d24c6b5ad29b0957fc33570895c2d956fb3",
      x"c9322ad88c5820ca4e7100d2bf838989d745910ab3fbd4a5b2dd5e6d95fb3c80",
      x"3156787697e9c0dde72374187f9bf5d69393a414bf5c38bfee3afa71b2982639",
      x"6e1eb2c9aa0ff371c542e061e4257a4aab8295001094b4b8c5ca06114e18ca76",
      x"adf2e14f5d132b5b93d1e2279db05b7b7a835b0621703ce7d13c8c02cfa5f8e0",
      x"119307e29ea4134b48c3d132052c6a60a47c27395fa67a8e9b26e04767826063",
      x"1b753c5b1dc63c80d72940a9169f42cb3e2bf98d39c9ec40ac700a5dc9c4885b",
      x"32951059a6c1d2d4d9e3ac852477f832846de7b3749e0d2615fca6075dc931c3",
      x"d64a72ecc017de3ec628b679a6f72b7552e3510f1939d36f1f58e1fdcdcfc1a2",
      x"1672c28f0e6b07664d99b7db01bfa431c002fe4cea1daa2f458f3c1c9b420c09",
      x"07565903dc2430eaad182e9ffa6d37528b5e47301597ea420b9977e51598d6a6",
      x"93698d8143174a3a255235b5f063a41006f1b2fb26b35a8a4b92747ff8b74109",
      x"2924bfc98c17d795075fb107593b0470240456a0633ed368649e94c13d2a5579",
      x"2d43cd30e1c76dba86bfdfe46e06592a8baa8f3002b9c79f217d91470d88e196",
      x"3ab9e5c2a181d908da1a7e0259ea9c09e95c0151096e43560179e03cbc2a58b9",
      x"2ca1c4e266b354502ce3ce46c6f5aa71fb486b513b3648a2c48ea57ce0d2a1c3",
      x"cae2df4e951a427270c4dd449ca69ff6c7401de8b85d82fee7de530a3033843d",
      x"39c6d2a1d5eb0c37f143e0c5547c199863de22699dca096f8e805cb7169a3c5c",
      x"8e59006ab89c8478400061db60cf0ae6b4ba90c5b2ee747ad6a76dcf3f33f576",
      x"3c970501b53d68a373c609ae81402ef7c2e5742861894f15a5436ae91a052daa",
      x"14345ea323a4644e272f2c70b723006506beaaada948ef03ce16366517ac47b5",
      x"a1f6f707f5a9e857657fd5b29b99195c77c0eb7c94df75f2e4808a7bbb23959b",
      x"59e0c3c0e4f44e70003444c2e9b413c35fc084075d6a957bddc0a0882fbd517e",
      x"ea60cff0069a90cd7c8aefd0bb9ad37558fb04716f5ab609a2202e4f564c8044",
      x"e5b012e8497a6345dc6b1283e49a9f1e7adcc12c96786f76d972e2fed7c40dbc",
      x"7914aafcbdc1a2dd28ead4c858756e619899bbed0c15b3959dfb531a3256924e",
      x"92f5651fc28fa3b7e2b8fcc458a7406c4f2f83c4ba7a11bda869da8f9f341698",
      x"9b0e29978f02b38d4e4a254c625b00ec36ee3d2a43411761efa335a862df1ffb",
      x"8f5ea62e32bf65999e83e87151d11641b9cb9bf387dc66501a2166aff27cd40b",
      x"c57710bae82ae7b14fe90a96e2b542bcab5b2500a05daeab2846f7a1ae577865",
      x"b98d2f8eed17abf9fd6e44183f913c2b1fec31176c5b9656864709bef2160f39",
      x"07ebbc9b077242e25330eb1dcd427a99b842fea3fae21f627011c1c8696459b7",
      x"3950f08b9e94a5d16b18afa0443b38fea8aa5caffd2d5bc7a86b03f24c974047",
      x"9c1383f237da9d258bdb4488a861b5091e78ae282fdf2586a1554a42289162b8",
      x"f89980fb7c91c9ee2573adc41b6523373516a7be25ddf1f33a969549cf5b9b09",
      x"1a9481e80134c4abfe4e96757aece7fffb0c5a3b2c33f916ecd19ea344b0734c",
      x"627121a053c22302b4bf026b296483d2f416f3076de3a466ebc83195fb0079fb",
      x"05ae4d19a9b51ac3ee6bbecc7079b9b93da505bbccc28c36ba3a23ca15abe276",
      x"d0b620b9d3140c784655b929fd8a2afbc52a2d4327bd439c34399776c6016b3c",
      x"750827a5b28bc0aa1097a8855b91847099857f468abe2a914e335ea0323cb502",
      x"0d0d2bee23a0abc557d9b028a9daf77059fa8d9e8b5a167038f1cf2b98893d00",
      x"ac131f8f41caec2166f3297ba091e227e9f06ad6d64ba1fa28ba1e51b1e5030f",
      x"1be5269a0e36c227cbcc64f68fb32c3818e38528fc6dd8a20ff56937d87b59b1",
      x"2b5a159eaf9a7a2cd38f0bbd407a14dee23893f6f0aec2f2e091aef91df9131a",
      x"c3c50d5f1bbb793c209f96d6b89dcb6e7963138765735b42117c56f271785f5d",
      x"44114b982276a5d8001dfd5b3d8ebc89121be15857e464262bd4c51541017b85",
      x"527b55013573645cc3bd3584e2f1246f96f15910b5e64478971bbeb73752ec4a",
      x"51680d72110a9e9daa5840d49affd3d90908cc1d60e1118cba2f6b48f9fc776e",
      x"5dbb787676e85b92c08d0fec709f9afdb745d6bd7ac0c4237e35e69f5487962a",
      x"40f6df757806ae4c87fb4ad38159c50ad44992c4dfc375a262e67ae495aeb1fd",
      x"badd76ea68b57b1a38c710c1988fac98db53bcae5a5d0880ee5149a98a95ecbe",
      x"bca220a6c80e4aa821e3443357f1cd4ee2bcb59bb7933cfa739f053c5726bcc5",
      x"e7e333f9d648aabbeacd1318fe7eeb41313cfbf000d956f40455216d9e444874",
      x"7d5ede3fcf0f24cd65e8f440ee27c2246d76248921f15f1a7e6df9a9eb7c5705",
      x"0d03aa2a146dba59272acc6f56131bbfaf29bbd9b0b8a3c6330f62ba5e94d24e",
      x"dc25e8968ea468543620326017dd5beaac22b34d7ebe4a3d956c442aa4d5c662",
      x"c14306d42db7580a2f54164702e6e0bec2d770b4c17d7850e1ef7a9e042b8b58",
      x"00ed2a5597c18387246c02d80390d0b52a855cf42e3c14d4dd0332b7e7c150f7",
      x"ebc65f88a2ca0943b403ed0e8b96c3f82e9ee574643beaee7d9e97f9d683210c",
      x"c787ad4132954c5d52e19e13c6db384b18fbbe6d51c991990b744976c86c1314",
      x"f38705cff88654012e1523a2eaeb60bb4d29b6156fcb8d5780c5ad716b8a552f",
      x"1d458badf3c96a6b33c309d98a16f8247f6e5cd8283234b1e6eb8d8c7eda6510",
      x"aefe63298542db59fad8c70e4b8a1e3e53b721b30bcea6a0196fa2ed0b53dca5",
      x"cf8d9243b7fab9b3c3cf5297f84bbf898630f2299d07b0fe09a6be2a9c5fee0b",
      x"6953643a8f8059fd68991e519972f4aa3d480ba6622c3dca2fca3bea596dd540",
      x"1c65ac418e054bc9e7c2434e035b3a59759e7f1545ff806badbd1208a8c70096",
      x"9099d238f8b033ff2763d5ec17e30c1facf4cdcdeb647fdbff7afe72c9c9c0c1",
      x"5265501b8cd2275dd728bea0ff638a5fdf2dd81b997ac53473323d42e3b43276",
      x"c2aa77cdf8ad98b73647cbe676fda5ce9285c99e0a5b2d3ec330c56d7e74528a",
      x"df483f918331379b14404417bfae7182c82723d8a697fc714086258d1668a8cb",
      x"cda312c3f5acd7e195e132fb75c27f2fcda4069069fd5a83b9bbfe81be710e38",
      x"c4becd9907685744d089a6ea4ab1a35035c7f885841a3cdad1ff90323bcc9255",
      x"15c146c1dc9d534a98dfca1a608715fb48a56284f265aa62b43b2ec962cfaf6c",
      x"04ae1712e6b34d5393ae0463b6571a3f4498b5fc84d7ff75e5d10fe51ea3bf5f",
      x"b0d592f35f3fbee9b58e70392e4ae467823c50e4b7d321f22d243f9bf4bc21f0",
      x"85cfe064caf4a28899212ba0b63870160a4aae446f1eae859905187072658c9d",
      x"7773c69eb3b54c6a8da5f1640148ac3c131e88ff96bb2b3a14925e0ccf4bb573",
      x"1db38ba802619b5a533a0b78f1a5cd5fee8ce5266b092d063e602a006354f482",
      x"359c4ba47683ab36b963632145e52ef2565a26c4b6121ef9ebc054b9994d4ca5",
      x"1b0fbeee20b1480f74dc1f07b56c4346af1c63885086b4c7131bd0e9fa7fb87d",
      x"ee5116e4832a5c23b30c4de1ced1abdb4fa16b224b017477fb61d6bf82ea4a35",
      x"bbba25e2932a57791b4650d151c76912ac50f246566b57212c171c73e7729114",
      x"77969f2dd3969c9622a12b52830ca06bb684a1ffcc53c5d4cdf52035719f519c",
      x"6fb3471485db9f579cb0bcaf491f31ed378e78e5d6007c41570de5212fbdf370",
      x"8003b81d886680bb14fbea334faa54238c6083de9750d164cd1e7656cc60a9f6",
      x"8a42db1ed3828fc12ff306dd67ccd6515f4150c0e1610b1e12a48bf2f4a108b1",
      x"05b582e9a88799dd7ba8cfcd405ae3c2511418edaee21701d7e9b04a260ad39a",
      x"edb5a6a39e6c74388ec793de68ba1cc3910529d049093843029058248273c498",
      x"686a90c42af5217999a0bce17a983ebb18dc532f8494c2f40c0ea9f205a5c620",
      x"3095964e526961698f657c3320d35491a3c72aac1b6b6763f457d27197d5575c",
      x"1ad392e9212dc56848a98ac6c9e68a9df69198384f397cfc1a13a8e029be89f7",
      x"7bdcd940803d41ad435aee5532728f978d483e2b5e53e6c87e9522e17b8ba631",
      x"ca3059af7b1a54fe549d2664e9dc288cb9ddcef9dfb711246bf5812b4f487f0a",
      x"6a9ab4a85ecbb13baf10c09c982c1a1e8aa2bca997e2f71b16d89c9108431db3",
      x"152201526d538208719bcd70c0b5ee1382b7deaf568a6cf95fd6a29d96c08e25",
      x"6a63879b00506504fbb4c27022c698a3dc1b253f3d6d80430f5f2e8d9fd15344",
      x"e805556218a2df427ec00b31ef6995a4a0bf4d8997a10438a2573d5363aeb33e",
      x"9236be5aef6830d68f34369b944fec144e96c9593626ba1b5e15a8055a5eed32",
      x"21ca32a5c8f7d9e0b85e3ee77f6acf9ba01b2ddb945ff7557f6dc9d97bd081ae",
      x"29870e4eb68d471320c4d9bd495221933af3185ca3a7718e8f253d3c403cac40",
      x"8b6e5b5f7fb41d81505f0c8b0abf8736bbc9111df030b59708de2db75cb77598",
      x"7b8be7a075652b049ee56c4fe86e565f1731a50a32c5f73ccf690c6324d66dd1",
      x"29ca0ebe38267b6e23782ed5fc9c23cae651e421c92a9b4668c3401d77c3129d",
      x"36f480e3b69b17f8d87dd60a83640f9d2944177c1ae77ef0019dce1b8840f576",
      x"30816673260a8d94e581d712270cfcf37573aa27f876cf16061487a7ca6b18b7",
      x"61daece9c76f0d113610f39e8da003f191ca347e2850db69f9fc8682dc61708b",
      x"af861911437aca4648d2110e2bacdd726988f2e70183078c44b2320d6e20726d",
      x"24e7a6dae85fc2b7a239b99891daab6a9a965ea9e3486b7af15aade22cf2fa7d",
      x"c0d004bb36e3d199d3a0e6c96055d809bf7a36c2e447d4cbc840ea2a5792f632",
      x"cadc57badfb40f3315bed5a2dcca3102f6a8b4346d270b6ad3c4999ee11d86ed",
      x"6b30480c6f3c1b1ed7c6523dc3b6c83c5c56a3ed7b70e55fc9967b89f4fb5d81",
      x"3fe6305d5310e69e4a77a20b5f8b5d0342c31041df445fbe084b92cd1e1f1985",
      x"41ce0b4c4b1d813d95e42c7df843724458254d66d2f651162d52872c4f9f3d2f",
      x"e6babcc129a650a62d23042ae0c3a4367bf0484852876dbd8ce447ed24ffd63f",
      x"dff2dfdc61b4519e5a987069f685d697fae897afbb990def8ae3996f82ec7f2d",
      x"a1bce53341d72b41e7a439fd2a13cb724c47b0b9a95b94bffcf59ed31c456746",
      x"ec67ace0eef3b55502c164065594faa4dada0f5d3ec07fa10de10104f4f4034c",
      x"45ac7df176e55cf3f4552f7b2395a1151d51b0d54481b8b87fad611f4097ead6",
      x"9779189368e66d4e05c64b3fbfc9434fc00f6808206a7564414ea33e6301b17e",
      x"442e4ae23440e11b316a3c62dbcf242d5236d76f02a55bdf665e51a445d0d2c1",
      x"8c3da9925e8aeec5181727f8b5969d234ee6b1261ef7a46dc09ea55c25018b7b",
      x"f718ef0b787dde5e0fba2f27b1554d1a45f4c316c4115cd0b18ea1f91efeccc3",
      x"15dfaf7e6e0b8532c86240d9f1e99e948f1adc6f9b2809d59121900278c97ab8",
      x"0760d1f8102dc5d0399c7a17ee387d93ab3b1da26fc957d33c32c29e35a299f8",
      x"5c5f641b82d81c03b41d9942afd06cdebbcace0e94e40428a79287d8cb438c3d",
      x"5b716b489665be4c27dcd246dad69a891b0962921908d512397b7a09e5214341",
      x"19acd43412864b6b2a99bc4eeadcf76427b4ae01f1d79673d29317403e5c3273",
      x"0fe2a2a288e60aae1f91e70612100623b484f8b9612925baff83063d44ff9438",
      x"6507d0493500c6187fb134fc540d6666c496cfa272e7558ae2260ce749916f32",
      x"064ba13de52720ac41444cf832a1706ba86edb8c935d54d350b849055edc77a5",
      x"3e9c972cf183cde3b2005fd22cfe800f5118ad412821fd9d87def747c478d9c7",
      x"c55f71f528ec3b3df6a6a7cb5bf42e2db2b8305989ebacc9ca06132de9d24e9e",
      x"d97e3d7380ce920eab4a57f2ce89d53e55142e4f958e4f85702bd900ba600ec1",
      x"78ed6d178a5af497c876d884b52309422b56f07617c72a3c0c486511c7f05c80",
      x"8b52dd9dae3996e306523be18d6a0d4a2f69edc633bdd65ab0ae27f3aeab21a8",
      x"32325d83066522c1252b4450bdffdae2a68df9485f3b01a1ca723aec8d10da5d",
      x"47e06ba1192417732898085657ccd5c9898b934a3e09c66216d5655d48d2863a",
      x"10fdc00268bc3e57a1d55a216a4bd49df260637cf28ec79a0cfb8e3d15f0d35e",
      x"2f8a7556d48d49b98fa0ee2104d8c4f0e9ab3a5cd5811870bfcee7d26b9dd8cf",
      x"7d1f9b2c4b4aca4dda627d5cb8fcb44f990f4122126357e0e1d8c6135e6417ef",
      x"bb8214fa243aee8318a9523018046b4c6895bce14809f5383bf203e7d62b8557",
      x"569aa92294b2116d016f46e69879b58f9cf48fd29ded9835c5e4f20638040a21",
      x"ef660b366b15ed717f8144cc7915e6d36bc6d36befcbaee735407e57f8a5ce02",
      x"f1a0fe65d755b35d297eec9041efd7ab524a6bc30cea769eb45eef2b960c40ea",
      x"e80528de4a245ff61c38e0291b6ec460e490d7a4f6a796be6cb93d52e5af78b2",
      x"1f86095c4b353a6fab09fe49953eded37e6ff884b268978adeebb0058ec6bae8",
      x"d19aeb504922bb6a845e12883ab38de218dd66c9485039b480a2654125980cf6",
      x"09dd5e07b44c434e39986fa793825dca6c0fdcf7d45ca9a0613203f8252edfa1",
      x"d6c16499f2a9d1dd15db853a36c199cb24eb479801fae49bbe0669d418a75e8c",
      x"ab0c5025df28d8b32f4a5dc11cc500be5aa11cfbdfbd84a77160230d308a097e",
      x"d37b64924f77aae0d12a1e16261ba1efca92806f8ba8eaed00b0840e08449ace",
      x"5dd3f6b2e52ff4a5937cce462bb6e32c537dcd2f2fa7732c18914f192b3bd016",
      x"034347844ca65e5c6c5be5ae6f356befd480e24dc833eb7642df49069460a213",
      x"ead01ae960abf61a1888ad9fa082c57c65dab3c4db0f6cb1cd41226b30bb4010",
      x"c1d1bb00ac0a8145169c8dabfc8827e5e63a0f8a378beb6c65a42cba8f355f5a",
      x"f4a596a51cebce9d612958ab4b737dd1a517cb6b628ebf96f92f4c74bf1d73a2",
      x"d7f79e98fd1ba725433796cf34196cad91430e69a25226fab6daa62033488cae",
      x"ce73a0140adc556ccb550ad6d593c2a520ba9af34ab00442c2cfc23abd17b02c",
      x"8dc925e39db8b28ccdc1fbc599151b9d427738eb0a56260a7b43ef5ce51a2834",
      x"fb330355b5cf330af06676ab82988d81c269a1a24266e6ec75ec99b22004b797",
      x"f627050d680845fae6039c293e89e97f10170dd4558a71dde1b7258d2f4daf5a",
      x"6a0a4035d70f87252b376c85bd664aafa01b034580bf62eb6dd53bcad8f45206",
      x"bf4f60339e47d5c44b86c535508df875c5422ad2ff46563e1f163e99472938ae",
      x"a287891bd642d63f39662add8036d1054abbced53a4b40e002e5a4848cf18449",
      x"4179cd31fb96d234e4e918e370b1e4317fddae800afbfe65cce449a5a15b67a7",
      x"3421f0d066485d5878622b4002d7ff84404dfe4e3e869f0eac34eee477b9249e",
      x"72dcb1011605cf40ebae0a9259133f4a81ac9dc0ccde4f037cbe9a14f12e22ee",
      x"f36677061ca79e114caca2b36d1ff9b58c521906cc6cc37937b4f13d0f1e4fc8",
      x"4340b84d2e770ef96afdfacfc6ace4afaa150e368fe4ab82fe51d4f5285ac153",
      x"72db244fa6a0a950843e26ce5ef7586965b74734744d3d36039139dde7f64e4a",
      x"0b6e616e9072a1a0c5814ab5406f00b9ffba042ab5844b2d2d605187a564bac1",
      x"0aba93def581cc55791cb616ad4af9d5ac682b07b205d9988dfaa0db2f27a2fd",
      x"73eee7aebf34b3037116dcbe39e1189e9840335f7e1f7145928c0d523b7b0544",
      x"4eb7bfdd3a4b91c709134a79f429cb4ad361af55993ed9ea76d41b9ca57c30d8",
      x"3b0ee04de18badc01ad03ba84d4102ba5b35ad5048f148bb2d25165f42468093",
      x"3f84118441f660df36ce4076049740f19d10dd469c656a611fb23c0f81159105",
      x"215c0c8bd2ce33d9ce97df3e3d575753db8f0306e536a9b5c1c3c16afd28cd6e",
      x"03f8ea3c3e334b56dd762bf5007bfd9a5ac116e9ba6ac54abb295dd5ccaeee2b",
      x"f12107d61f1205cb2e02483b63f62bfe5fd8207aec843e4da544b907dd9ec343",
      x"4672a706dce027b2ce16f01f56dca7469b304201068dfd2a04b33efee93ff630"
    ),
    (
      x"e397e734cf99cd560cff1692b8eb4b107c43683df08a40ca206e632f05388823",
      x"cdf5a6a1bd75c108a44ba7e34ea74caa7369413a27b659f0f44eefb780bc13b6",
      x"54adff11233a60542934e2a374b84ef4c72a3cdb785e813f965c3b18cada6206",
      x"544b791d8c49bab29b7640e9f12cf9851a33d68404883ca27888621f676a4b5f",
      x"3524ef2ce14935f8d2b3c403f5f23c34089cd40dd2f028c838c1e9af0a6ee9af",
      x"a74610a3de4c25ad2d13a407bdd205592e62968e16044c539c8835519ac1bc55",
      x"f120e02c17a1e8be9e8f90512d4b442994d48bd54a9ac85a08dd5f2ca5dc42bf",
      x"a36f0d34a4d8ab25b7c24a8ab4930236d2e877846c7d47072fadef047743daf1",
      x"ecf97a39e3e111a31a98bcfe8f2ebceca132c457bc41cbbe8db1a92ef56204a5",
      x"d2bba329f2e02b266bca75f6df6d6e9864a5f57d04e5d0bbddf401e23c25acfe",
      x"32976ac1760fca17acd671a49b85467dff91eee3353b9e66387ebded2a07e5b5",
      x"1360f9aebd5c501b8e4edf9d868e783a2ca9624c8e463d48a7f7e4fb857b9714",
      x"bdd07cf5d92fe71249c0ee2ca5da1a8cb8d0d82cdb2e98353a3e74c3e21611ae",
      x"6c923fe70bc20c3daa03bf4bf9455b9981a659c6cdfba1e8d0f4f099f8b750b1",
      x"cf067a9de4492c31e284906cf7ac9ef6f79628ab2a41166a1e11073e614b5c4a",
      x"3cda51d59c608c7d287fbf8bbb7299b2153709fc72f6f17e92a212d4a06a0b20",
      x"94f408c33c5ccca721a2217b7032faaea4f6ebf8f0d1ae12dc174383f0cddcc6",
      x"cfed45f7985b7f8e1a2a13355df74385322d30f84d2bada9eb265d3bd1ff5716",
      x"8e8a3372e7463fe8c8d82c0681be75e1ece1af9017a555c9a031c533ea1d8f14",
      x"c16223c9ce1631fda77b6ca6dd5d3942496feee651699293db26a80dfaaf85a7",
      x"5b1ad79a0b4c0a4f8846b4c1fd7558256ef26f1f15ace9a704350069328a325a",
      x"198867a766af098018ae8ad064991c2d52ed0e89ee8f85dd17deae8b4bf914e1",
      x"54a18dbc8256ad106abf971aea7c833f782ed6168be8003bc517f48cd0bff72a",
      x"dd1b52ff397034eb304630e742e4615f62d4c3ea3d7d9af44a9c96d744ebb705",
      x"cd3af1302b63d179daabd066325bb0c1001a2a17ddf052908656fb48182013ca",
      x"1b4683f05d6d10299b0d5d5b7de6b192be1badd776a895ebe817cb01b100565d",
      x"91e050adef65046f39becf46b52c72f095cfc5a3548e070c936a3c0fc738199d",
      x"66f3680a44c88a13fd929dc8508d216b9a7619991760ef88182ef015fc051ebd",
      x"dc27537ea23cac6903dfb2d97e2064fda0bbf4426c5e1d1fd1757a14917ad8db",
      x"9e3a42a210548d32c8dd2771f0240073fd5190d384e79d25db93db2364a0faf3",
      x"52e5e72a56547dd4a421122d52d5daa9d9d41abb49abb63b1a58a8f11cba3837",
      x"76dfafad54615eda1b24b22c5917ce2ae4139afadad5c45a0571f9f38584dd46",
      x"c4d85dbd1a17fc27f929de1097764262619240ff3ed8894e74a55361a44792cb",
      x"2321f69f52d00c7e1f0b646790aaba7baa26110c2bc6d4cf5a5eee54cdd908cf",
      x"157b49d641a8bc82aa3c54bb90ad0d8d5995dbe076d151585c60b7ec0b8dbd9c",
      x"d35e1377ffa8658027b20a69e1ad7b8e88d9ce92e97981a4f34261c08b589aeb",
      x"3a083119cc47c77e2d915f15891f9f93a196d9342dac1a8b9751f4c91a34b17b",
      x"afe5f5178e60cd0efba51114eea768a54c72b3fb723489986b708f21d709d492",
      x"a992536d9ab1608a8013b81d081bc4f45e7e3b38055359394cdc6f12f148d3ae",
      x"68fcc3e04689da2b349f1818707ba5a9b6799a713f2daef751b381d9f629f8c1",
      x"12619be4aa3a6a900bd27b352088cff7a7a3eebdbe95455220a1e8b9324b5166",
      x"554bb80812a1d17065a3a93839c0b9b63150e2c956846e31a448930a0d0416eb",
      x"15becb1ab689c20c9d42e8b7aca07e0f4d9dcf89c090763b14bf60974b0cb312",
      x"0bb64600f210f4ccc1c22542e0769a4a0e40628758ad53efc02e8aa3e1472d35",
      x"25b3864cdf3c9072f49eb499620da3b14e56ab2cfd0ae31469560dcf024499fc",
      x"cd8bc5a1cbcc20a3e7d5170e998ae0255d3a334cde7c37cf2a4371675a3e4d3e",
      x"05cbb75a82e4ce20ab574985bd425d2a73dbae27704db2a423065bdc22a7abee",
      x"9e647687aecf2c7752f02faa748e9a7506ed1de0969ac1e6d8171017284c43ca",
      x"0fd56c3d1be352b2199ecb9cef7877f90338bc66bb1c735603bfcb6766d2c716",
      x"37517eee933c614256f96fa141d7e1f850df757ac8f58c221383efaf991bec7f",
      x"ae6b5ef245f9bf038159dc5d0e148ff9c665773247ce79fcf0751bdd10cea8af",
      x"0a9438b09234ecb3da61050936b78f76eeb8c1568f66d10ad88130275d660cb2",
      x"f6543b070c2b1e49eee12e20366bfb0505e310b46ced2d129aebd94d2ed9d68c",
      x"a42e2a6efef4636d46d2933ea93750a8045f69c1cd78847235447fec1bac4c5a",
      x"e6fac71c3d56befec3d2179088af160d72812c8c82b3b376d611e5c9f278a7ca",
      x"1f169322da3414b9ace2e4ae97136308f8d0600cd48f5bcabe93cf4cddc4c58e",
      x"6d124250c38bb4ae4ceed743fff3a39b417f3eae35b0f1c63cdae7c20cb9d805",
      x"3bc89cf553132fd534316773da9b82552e04e7cb8868d8cac6056bb77df0d886",
      x"f15add833a4f5eaffc67e027021727536884b05303e579ec51e6762a5a7b2ff0",
      x"f9963b1c6d0ad5102bbd32eef102460dd641737ac6ab4922b90f3d4533dea126",
      x"e10593f05a5785c20a92192c60a44df81773c2ffc410f2a3be7c0570c0461e33",
      x"50ad8542669c9ff9f521d33a612f6f0baa5e6eba3d2c7ae004f91b31d849f1f3",
      x"513fec30c50fa1d5bfb962b6a64313325b6ba180f2a9a6cfc3b76f791914a78a",
      x"4bf5d24607bb59b7492dc7ad86e83f2017fecb2d7f0220a4ff38ae22544e2f55",
      x"03d0783a9b37f225d8adc44c559b07b0f5538c202054d29ef535813d7772838c",
      x"e692099002c7b1703fa01d37106b016c722b43a26052f685e4a1c15bf357ab2b",
      x"ce1bf547a626dea3e24da1c0c08566811780466e0c8045b52a15b313629de8b6",
      x"e1c639cf57bbb79ab7a65be4e177c6242c11f781ff5760c1066598d4736178c0",
      x"6984a562f62605c1b1a5163e6ab515363cac77838b924cc497777ea7e4c40d2e",
      x"55c75c94fd873fafd84e678922815a230abbd7b81700ba746d8667944844f206",
      x"0bc5e60a8a6dea45c03b6f26801f164f80fcd784de0037b54a31310886fe657b",
      x"bb495ded3a78f7bd3a30a1ff9c84a039804fcb72336f5abba9457229381dba83",
      x"0949c4ee0f6131c1c511291796cc585a53c96896dc09c3b3b1ab3017aa30e431",
      x"3f48c63349b1168ec3de738ef0fc864b383da1535cc9999970f3cce7a5d58b5a",
      x"ee3f70a31b544689cd89cabeefcbbbb89693ff7db841a90bcfae24ad6cd1e65b",
      x"21d53904929ba6cf019fc6c8e5d87ac2e585897718b0b18237b3425e7fa84e09",
      x"78a9ca038f1a8debc80f5b8d2ded5be800b8d05cb24707c333a46c569f8c6011",
      x"1f8386a81c77aaf072677b230baf1d912fcca2297606bb71ad9e207cbefde355",
      x"97a33f875a0ac2ca6bcd3d14ecd1d06b0df3517caaaea544e1aa2cf13d8672c2",
      x"35486499f5c62892e530f749c530783eef02a2a0aef8212b87c3ff35fc08399c",
      x"a9edfd2ff4c991ca08e63c43369135674077b7997c225bef25e108377606a8e1",
      x"2291273a901ffb71442a48b9bc2601007dfc33986dd3fac6747f48a6b7ad7e04",
      x"6c914808b53af444713665d383710334bc0b3a15e935f8d3a2b65f31fa3a9633",
      x"945f719500839bc8d0c244645c2348c0accb29bfa602b60362bc6389d875d9b8",
      x"64295fc18b9140ba10abff1227f660e5e62c8d75086d26d4b16f0bf3d1848522",
      x"a45bd9b1f33d35c5ababd7aa20276a5e8db2f176d18b0e9fc8a388423f1b1db7",
      x"e6fea7734adb2be3a4a332851e241d5d0422b97acf6d33705f398336239112f7",
      x"0085cb36887a613d9021e317948635d145f1cb3ea550483b8b7e5dec9c0480d8",
      x"bb070583bb208b776dfff3a0cba60a34ae62ea6408104896762d3a74b9f0d3cd",
      x"ebf207ad90a47e9e38bdbf0ff44521704395ff80788d0470a83707b2b04610bf",
      x"1a788797dd1f349f1dc23cf85b6f825aee3d1b93a65fedfbf638c5364abaac88",
      x"c0cbaff55aa7a6c83be4497ef36393bbf741f26af131ec2f4bb3f77e6cbb8f49",
      x"c61660d7641e72f599d4560b57d6241fc54ab98fc7a3029a475cecc34fe5f2a0",
      x"dbbca295ecd911b43fc06b2201ea1649412288a1a8d73c1c36fa871e4a02a1f6",
      x"66502e3793dcac4e1fc39b54fdddb45a9eb73f460a2b99d71e71769f7bf44591",
      x"e527ac3a0134fae75021926fd54c1c56e949fdaca9226c6bec61a6b11ddd018a",
      x"870325edabd229c0f84c267904323d8ea9e8342b4e763bf64154ef5aa8a92354",
      x"544cef362f487f004bbde6fdf7fc63e4cb269d37d729c460819f1e4d09b09b99",
      x"815f114e6d0f134ab164a05cb43940b2929ce910dad6abc8bb40095adfe51fdc",
      x"366b60b5775567811e99b694bff09607e1397bcb5659e27466bcc1e243bd84ca",
      x"15cc951ee7b70a086aa3d4550c1f6917e47f72a291c40c329c35f2408fac7910",
      x"4c0932fc8281b7504138e2b0317e0e0b40511b5b9461cc7c36e53cbfccfb56be",
      x"674e99c1095dd0c760cd0ac7bbbe713b0a17b5f7cc2ad6c7028146160fe89cac",
      x"1fcd5338c151880763b2c4d0844cc72db9a2b2ca5723078c0b2c978da5845b63",
      x"c9c8e7abdc040b8d246d1006a1c77d45223a8e1415f46a9c3bb89a86716e5f6f",
      x"0212758ee596087becac0e6e4c251558b4ffabcdb40adaa009cddf78494565d5",
      x"b71dcbaf0fa49b7104c3b00b10f50661097eff78aeb0a24dd41b528f73150f44",
      x"b545a3ba05949241ac99fb6b6a76855baea1b7d14bc0cc635e44860cdf889278",
      x"5ec639ea1a20e214924d17eb3f3697adad69e5247904783fb895b3e46d485a1f",
      x"34a0423afcfa6a52916e610db172393ac689fc6efe699cb1e51b4be5c8afdc9d",
      x"e96b2afeffac4ce8f15c6c52030c17f9370619ef14b4501bcdec5169ac7b1400",
      x"8cfaa324facfa994f2260e2f099c4ce27b83389fd1f93f8dbe538c00578a5690",
      x"e39151654da44bccc040f5b9ff29e324c24757ecab55873d79f4514921de23ab",
      x"4bfd496cf4687f80fe7967fb1b510fc0d02392086733da78a1b7d416bc26a833",
      x"6c6fb47c2c22cb5ec009eb8983bc39b49f60eeee179f1172d08c98c47c185ae2",
      x"89fe54be9e092eb5d73d90ef14cdda1dbcbe9486c8e746beabd48e3b2d55f7bd",
      x"d3947df254c915695fcdd7d4bc0098ff651d866d6ef37800de6323038eb7ef54",
      x"2e06d89bc7e717ea904b7a44ba04b2e0f42e508653a1dfe59f7a997d50b61536",
      x"24b7b5193e10dbf5414abe37fcaf1e1e8593cddf71d07687fc3ecea082a8631e",
      x"bf864fd3a67d149636401996d4dd6f7bd7efefca362c0f2bd0b89bc1f07f15bc",
      x"86bc68a104552588695e50290f4a46572fe84e61a42c8ce345d1598e48208bae",
      x"c0dc89801cede55839009dc0cf335191067c8c50367e0b181609b424f3e39902",
      x"2694725047194c0c3df4c32d939c419864b4ec8492754f161e52e1888b7a9ed6",
      x"cccef2bca94a3e2ddb87abf7688b1fa0be0d63ae5bbff125d81c277c04bbbc41",
      x"7681c09b0a353eab7acca72b03242efd8d45b8d44a66f73ceb544485b4aaf534",
      x"2141913d31ffa6caabc4bc644c67ca5d72eea5897eecc51ee8b3059480ed6c46",
      x"9b289f4d085d5b88704bcabd9888d3e65cce6023bdbd61f7e691cabe738462db",
      x"57963dc23518e32e56cf149532132f634f1e03ab8a092f4263bebfa3a766b255",
      x"7a03dd79b69ae604de2b1caf7397022578ab7ca27b951e25537c3342def681af",
      x"5ae3eaa5cd6014ea6f71adb798dd8d5d2c7d386658f97500109ed9ed2edfe842",
      x"88e5cbbc87fa7f5880ca614eee0ad24b3b7cfa3ff3ef7d84bc87f4c8e97732f3",
      x"8f8f93452e7db60e8cdef5e3e7c0a4cfe4b52beab20392458c7784a569068e83",
      x"e9b7f5fdae56cd4da550f52bc73177aa2385ad566fce2441683b755e671e4330",
      x"bf18a91f3c53c3b80b1d9f471b55e042e2197df10d117a21ae18d88989ee3a22",
      x"39312a0aad0e53062d5a6149d2216212e325e66547e2c19862648eb775a1e302",
      x"3ffce807fe13a7967a17144d11cbc2e08f240459b22d65ccac22ef054fb11d95",
      x"7644a05862708f818c365c0641aaa16b0b54f4a589689d78c87b583d60ee8623",
      x"87d70cd156104c3b07ff742f6de8ceef7938cc5b5a1d9d0fd991b1ae6db8c549",
      x"77a99a8a7b04ef1b9675970bafcef547e22a8122a7cbd3b6982e249738a5e67c",
      x"92fa4ce9fa8a0dcf3e450791b9b63b6aed22c05e934d23a7163bf7cbebef224e",
      x"dfc135dcaf20e706a06788f5666685d98d016daa636d79eb549fe0cdc2f63147",
      x"3d06646c57220d0a6eb8b4dcfab4de83c710dd2a7743c3c16aadcf31d790f0ae",
      x"57659c65f386de774da27ef8a83c5e562062f187bb7fa0a6f7f39627c011b275",
      x"d74219e3fea519db499ef296dad3178d98f1d1bed483de66ca86d58fdbdb633e",
      x"c5f98792c3a8f458b048d79232533de7bfb2fff1f88824bb3f1875f2eb7309ca",
      x"eb8fe90364d3ca548b6abb92d84104465ff8cf156a720dfe953d753ed1d119db",
      x"ada18519c865b635146e9cdb81403810647ef0cd5571529b39a4958a42b241a4",
      x"77da8039c681ca37affa20a2ba9d11de36fbd762cd96524b6f428e181c990619",
      x"5bc813f2ec11261ee535056296e5f4a6094569f85f3918be6a413ba70892bc6c",
      x"73437fa05447146d87a15a41c6de08b0108e0ce822d88fcf405372e37a9d7b95",
      x"c4853e6bd062bf75b97c31351d7c815121928ba67b08bc7b68bffefb1cf91388",
      x"40a0f94ab4bd598c017f80921771ea3defee3ed98ae4d4f3dc049570b2a250e9",
      x"a6d15df3b6a75c221119aa73d628c269a560aeab5372721143581c45f2840b2a",
      x"b64994cb41eda004427d21c1190aa9dc9061cb9a6fd937f2ef420f55190c7551",
      x"7240c7ba23d13123279c0459d7ebc5d907ade52e11a1f53c3190b1164f9d2def",
      x"59ab1b5aff003fd79e4154d36d51ba2e65b722e5dd551308bbd65b8ea14a31f6",
      x"621afa74eef6db62be48084a15c6c182ccbc95441c7e3ff8ae6060c7594f08b0",
      x"c36a65b4a2c6f84278eeee3e1de7bbef9137c92a98cb3d3b301dc2fd36990531",
      x"ad0a5d9e8b2683040f97616bbd6f3dff1be47a1fdb2de164247bf6d934c7948e",
      x"f32b544d227297c86e45586bf12e2054bac3d35cd45f08e2a0c207e06a00ce36",
      x"feee1f393ac346a64ca5cf78bd7702e93f81ca0d95cc84a7852aa9dccb9c7a65",
      x"f1b1c873a6093c2909312c721d515e496c3725f4e8a6a59f9870c84f669520f3",
      x"43d299609a3ce971f047deee59618b72848fcd5da9e55eb5754e67c94b5d5c9c",
      x"a41accf5ac00ebcfb365b4116984bc3795b0d6aa7421d13a601777a08591b198",
      x"210e6a1652c028d477d106ef5128f2f09bcef0cc77bc2a57ba50c891bab18fff",
      x"8d33c461cc186124fa3160540a15da51328fa769a2d6f0567b7b51a00abdc677",
      x"6791b3c380078bfc296af0c8ee8825f22d249f82e3cf0a058f7055bae09cf3c6",
      x"5e4a8aad64e06bebecb65dde2b22dbc6307cfdea909f9f967ef4dcb23a0e7cde",
      x"01f563fb0e0488edcfecb4367f16738fd2568cf028496699d1568d28cc6a288b",
      x"a1b23f1aae63562caa30094371fbc1f63fa8988bc6ae2ac3572dc8523b8c39cd",
      x"eb6942ff3d8edf0ea5952c42be3b56da88b8cf3f03e1fdd7e5167f2f26e3c425",
      x"28c0136110e07928ce8e4e9a207959bb03dd342ff39e347929f5f2bb54fb9ba7",
      x"581ae9e94522099e4fdea8a63f5a361716e77f3fd8e88cedcd117d5267daab42",
      x"86c13e2a86270387267275dfdb99cfdc08744e59a40f7f51a3153d8c35a1e3d3",
      x"8b91e47185be02d93afc26b6791c614a8d17e0c46dd72921e3c675d35eba3190",
      x"dbec25dc04fe39afd35e91c98671c8d0a8a77de7614558ec8971317f110e6bbe",
      x"646a8703826a1fbe07c7f35fcd3613f8586e930f71b155dfaae2274c53e5a147",
      x"232ccd9c3576f071a8840c7e4a17da221b8a53904a94e36ab61823cb99f2a37f",
      x"fb281ff72b864e7feea74d35f57f871dff1cf482198936161c5be298a7bd1696",
      x"90705dbee8558747ae8d1f5813a5a58f4250ce2cb5f75462890425656ccddfc2",
      x"89cbc8fba1e44d90dc28ffaf4867d4003e2aa7c6c0acaeb2ad64528b957d06b9",
      x"e862248f13979e45b3f9fc1ca4d58ca378de2db09b0a552912185c7ef8067735",
      x"25825585d94cc78e2afcaf06afc388d83c16baa6d3ccacc68c7cd409642deba8",
      x"29fdc9522d986a945b96250faae994a67427f7f9b8b780a9e6d8974a1280003d",
      x"c2ff6f70572135c34a8ab8bcc23dfba7db2321ea3c0ed6c7ec000028c0f077ad",
      x"2bbce148e9b17f19c1f5158bbc624108184511f5ca093ccd917434e62e7e2aff",
      x"b74509d42ca9ded1cad36234ad9ce95763387dee0d641e6deb62e7957877c56b",
      x"b3d1e86ee416d0854d477caaff79840fb0dac2c4c5a5b4d0c7fcdefdf7b4739a",
      x"49636a3f8c45c335d8dd698d2e33d69c2eef49e07b1a2ec1f35ff685e745bee2",
      x"01b224f49653e7176a7ce13b250a44fdbadf356184660c8208539acd814140f3",
      x"8d56ff77fc93443757e9b3ead8384c2c10355d3893524d3e0b3ba7c71db208dc",
      x"20730ea493d3216bc243c01da954dd7a3a01f4d922fdea7702c5e19c4c82b06f",
      x"9b099441fab4104b59de774719b4cbf7e13912fd48304a03878595cda5d21e94",
      x"c6225f87b7df8992f001b33ed1be386190fe1e6622623188b1433cc384ee35a0",
      x"28e4931f4b0b9201d80946eb0927619ca6041c30df11c011fe0e6fea8c7920c2",
      x"2480444a8946256f4cf7e1aaf3781d63830286f2a4fdb91ca90613c9a867a567",
      x"066823e5df5e7a5f25eb42391108d24da61d087c42fff8a29a25eead3d05fbc3",
      x"ba9eb72b92e6e9d2b8a86e99d2b00bf6e101472313a4d2a10bd3b822245844a2",
      x"5e697176cb4359eb44c115320b906ff33f9b48f37be405ff626e2e85087fe95c",
      x"22a46c6f5f95175c35110300a50d08be3599c542799ca8ee0091fc50ea6191cf",
      x"a76e8dcf107a8f33487dc9d84bd7f6850caaebb7a7d8159a06de7172b34df20d",
      x"a15a10c70940b04342bc18a46f7fc7c38e7ae02b3f09bcfdade5dfd9340171aa",
      x"cccbc81e189dbe908e65dce2d2b81c5d5014caca476cd621b655dbdac9e14f48",
      x"8f77f9d5473b2f22036e68a729e3b22985c0ef2507664c19a77a619af61963f0",
      x"45110db7898fc359bf7d7bd3bf5e2c4898bf56f4d8e585793623c47aa47e0e0b",
      x"ffa3e377510b16e8b9cee4a2c818975de50baf0617dc37dab21020671f0e2ebb",
      x"c9a876f0cc41756d7d2a1d60188ab65302ba7448a0a46c240a85f562cb0a99dc",
      x"d446cf33e8c0536a6dc28f772f6fc333857aeb296efba0b07f254bb12250c16b",
      x"bcbfde4049ef8b480784cc275bbd0868d86832fc855b01fc65e68ada4fc47e7d",
      x"36b59480d946844e9f7f026b43dd0578b148c8d3bbc406d149d2feca6167e063",
      x"b6b5f3cd4352b89c4378398ff4dd83969382d76e496f63a921a6834300045660",
      x"b2d20d4d72b86e2540f95177334a6d4050afc334eb6720b99ab15997ef55c25e",
      x"8b29fe487dc93af7dc33803a89c79a1c733eb8aabeb903c6d01f307946debe4e",
      x"82a23a4d004da91aa2efe8cdb5dc689876260c40cdcad0f2528feae05fc022c3",
      x"f8b7975c85ce12c8f8a501191b6ddd1629942c4bcab8d4ab0da18d41bac54a96",
      x"ae1627f66c7c480dbc3aa5983ff74d84471c5bac077a0a0efe9e868cd5a2a135",
      x"e7b1706d6ae85f268d4056399d4a83d697940f883295bdd451cd1c7a654d9c22",
      x"d3fb9ca6f3cd74cfc1a5959a1fa9fc56247e852b08586236f33fb3bebdb72960",
      x"0ac085ab9a53c38a788910912ab2061f47fb5660335278ddc3898d20321c2822",
      x"c69a53d597b0d8ae7636a3ce624cfdf0f0dfef02ebdc1d932038004b9789c9f5",
      x"b4ea7c28711c39a203ea6a2ef91925ae00c2bd8d44ebd171aeab7634f5159534",
      x"247ac957689537878c7b41abd755c89c42693efe9b35c84e3dbc753ce6fe8abb",
      x"6c037fa5422d2f6c2e7c564a8e1be93c88d2f2ee547acfaf29edd7ee66b54d98",
      x"9241f5771686ca57aa592f13a4c2f0df6a17dd851903d58bc7793ce26221470f",
      x"306049c9b5f0c2b42359660bd123f4484f3c83a865a295205fd6348ffba2db07",
      x"1c8abf4c2171799543e63a08777abc89c330b64477c5d114b26df80527cb95c2",
      x"e3f4d168f97645d4e458f7c7c2b845478703ee82f68fd2e05cee6c3d3b345391",
      x"e75a8a046d87cc186d234d8dddc4b0683c71fd7b4cdda8b3f4fbd7a2a488ead8",
      x"549a755d619a1fe6e10aafb6abca81f886fadddbf3d72bcc50e1c851d972de60",
      x"d06f731776f6a7b7b0ceed7e2c79f8ac9ea84a9b1ab7aff4a392e79c2a1a06f0",
      x"28d1dcd5490c9e70fd965f79c961ad21678b8e8caf52b12f9270c93759e4a049",
      x"12f910bab6cd6ff9bfa08840803927df7ac26f39edfd0bcf08aa007861144ec2",
      x"c57d1503b9e9ee1416597b59ebed6e6e6ea13073a1b93e170200d5d24d6ed755",
      x"b7bdaf7c5ec7380728a2f55ff866c280a7b5a7a7029246317fdf7ede915be4fd",
      x"bd160233e58a80078f6bcd65565b4ed1d97a4e66dba078283d08761eb4265434",
      x"f7524737a3fbf1b829fa16d6baded9a0af431b766ceaff2414556cd5e4726d3d",
      x"fdadcb3403da1d1531a365fe14c9c521e13f1760ebfe7cbf56197cf11960b0b1",
      x"ea7a605cffb1c5108becaee1a227247f0b7be0304a0fad71796d22c04dfde32d",
      x"84fef999dfee178d3b9f612575fad67e45b0de3f8cfc49add7d9751f546c8356",
      x"45681deec81ae9f3b7c37731e38562a25fd61b12ae25b55b79c1cd4ac38b6ba2",
      x"6d6c84e9ac5875944ad42f7139aa5787f3cb194cfe24a268483b6af63c80894c",
      x"c75e83837f1e2945daa070463956e0dbeb9d6efd35fef58fceeb53e5590cd454",
      x"b1aed9bf6678ace492398e0da5bd4d1143a8fa637a7c2996bc20374b0745b8ec",
      x"99ad6a748cebfa3bb3fcd82cce312e2f99ba2b4a1981dd2ba6ddbec822bd5b9d",
      x"8c9f565588c2eab319f9d23679dcb592b3ef1db03a3c1c59a8b299777ddc161b",
      x"49ac88cce2480d4533c28b25ca756e747d0e92d2d0695408de90ca15c3c352a9",
      x"175cae4299d04d546e8f56287f9824b182b41aca032eadc209bab58b0695569b",
      x"6e07d5e7e00d7c3bfff460b167b8be39f9620924a818df0a1088b0e5fe67c73a",
      x"0521182b289c7fc78342ae32bd703714e386d3f6d63f78bf5a366028d6d26a8a",
      x"309f484bca6276a820572bc1aaec2e5b81721d397316be4e4f587b9e4f0ef69e",
      x"1219dae0bd63736a1f48c60fbef72b56731beaa671a377b053b2efe886badc53",
      x"6a2034e7c2bc9d15a229f2fb6f368d13d1cfc7efb5ed7a09475b97ad337ee2e6",
      x"cbfa8a6f84ba8f55e93c32a59d1575aabdfbdb2b36f63bd07b1ffbf7ec35cd9b",
      x"6fabf3c1a8f1f914424476eb39930b84f04b6722d0836d558a25a9f7920b0228",
      x"1152f143958376e245cc1195937c8d8526dc38c28b05001130a68aad75d32b08",
      x"ae846d57c4d661deae8a27575be18400434242effe8f88ec0a783037ea001810"
    ),
    (
      x"16ca0ba87e0a0f1b03967b546405d93326105c6bfeb87b9ee5df7a8d90cf9e94",
      x"322d7573356c9c8484e6ca1d272a08f4ff6b9d88612011e5c405682f25a98a6e",
      x"6260fcf0d8cb37d63f0397dd91a472d6f983294a32b79874cc51605c415ccba0",
      x"9040ddadd318fdf31ed9ec1afbe346d65a7a1e0dc98797245a05eb5be71b6660",
      x"670317972399e137ec70cdfa58be1da04dcbed14f08679915d2d11f459e367b0",
      x"d42b4d818bd1bfb6004da09f70335a12ff4a1ed77ebd93fbad7d9fdebc1c00cb",
      x"ab857d3c3055fd3d0413eaecc8ec3c23f4afb33df295745b1aa1ec3c094bff74",
      x"ad74c81c60e02d9fe645f9ea971f88b42d8e88d50d3a03a50fe75ba4ea2b8d97",
      x"0d4a650e18cc1cfbe9e79bbb24a96dd67f6108832dd9e78558418a011daa5561",
      x"a8115cb673e678e65a976876c7e4591714780cd06887124133702feb1ca01f34",
      x"cb6a6c3bc762c3a7e4b5189308c4473b23f1b5b0828195d1ffbdc40a2be08ba9",
      x"1490e1706d4f1e31090fd760876a6266339b21ee4bdf3d59d76f5a04fc9dff20",
      x"172f5bfda2b6c7870b3753bdf2c105f161b4c0a3417e91804de4e5cb5bc2e326",
      x"624cbfccafff7fe6145fe698387c75867fdba48c565c3cf89d44bbf4ba466d0b",
      x"3b69d15dbabea93c9bee0733bbf91d4373b2788cc9bca082a955f2abfd8d0454",
      x"1b82e6cdc66c1f4bfae77f68c399bde8bbef40a83bae0676e3eb5e2ed7cf156a",
      x"8e86c79ab3ea77d729c14614fddb32de1f0feac9804703873da058b5298b8193",
      x"8cddb9ed09bd1a88caa5ca04ea2850bfc2baee1d4f1343853462612319ed47ae",
      x"74be7974f5f7dc98a6431790eb10c4f81e790345ec30f418f0c3926235df1e23",
      x"9e35d80a8e8685caf267e3d3211d3fbd4cbf44a93bdedb6e0b4c2077fca627a3",
      x"5cb2d2bc77d4f6d021fd9f4763a09e0a2334577e895866749dc5c55084614cba",
      x"c9563ded39970daa63cbdd62601eb6454778075fe13d44738cdf9f4b0f6aa1fb",
      x"1ecbb0cf0c7fde3331210c69a22ab3e74f346adec01063162cd2b62039008065",
      x"5aab1bb2df90269bb0bf21d4c792007b97f73c989d8ba47c3670f7a9b21eda19",
      x"50043aaf0acad2334146efb28cebc9d7d8bffc1cadc42e20417c0cc26a1fe845",
      x"f9de13399666e0a4fd829f7a4aeccaedde9e4b37eb98efe7a1cc5020f36f40e1",
      x"115f324879b97d0e74ab3682435bd1318b3e5f77b9f700bac4c48b00df25f8a0",
      x"c86fb1ce3279c73ee9ee6b91b77acab499cdc1d508eeb1be6d0af45a7fcd1cde",
      x"7d811ab35eec617cbab9f94a4b145da287cdf73869e9a73e0a2ee4f4b9225a4c",
      x"64d9c625aed1cd77321a020a99b20051c7d4529a2a809cab1ef5b20627be88f1",
      x"7c09b84a5c0923142f08c31859c251edad3e718839b7996a8667effd427a6595",
      x"76f7f81bbfb126cc5d03fdd68950a9551c42daee5ebec620318c5d829afcd814",
      x"638c20786ada8c2699727005c2116bab0d0e3dfa0aba25cc3c0337fb72a55762",
      x"1499af9f107301484614b1358656cd533e7f6cb1c869a6eb2f9e0f118bceac7d",
      x"38f8cd0d6f803876d7fe83f9841cad166893d7a20234cdc72cfd017b531043b2",
      x"842a3a00e5978c423a96983d83189e4a60746ccc4add39fb203097fea8ef7fd8",
      x"7c7409a3bdd2e8d534bd23ae6585b4a751f485d2368ec169de38e300b14b3a73",
      x"4de2f9c2f058ef9c09f9ad42f7726aec6039eeb7b28837732bac90140811deaa",
      x"c5c49b75d82d80089a95d78ee4387c89f7294f0f89b3517eecfa342d28e50356",
      x"c151e6313b6260520bf1876400ce28ec882c943d8a3006112e65171906debafb",
      x"64c9e5bf600acdb8addaaee442bc2e6f55b6751663655f8e6a933e4447b2ad9c",
      x"c2b2ca3f6b63e7088bcf583e06259c1215c5c0f1bcc4ceec5120a994af9d5c0f",
      x"0106565e6425aa2449f6475860f87559e17feac30fe074400b699cfa5865e62a",
      x"fb65d5953198eeb32b6b355dadf047a527952363365f885e0052fd771de6d8f8",
      x"623d4553fe63fedec4b0e407a2b90a4d2360d3a0a63ac05d3c9f1f5b86682208",
      x"e6222d41a5fced62bf70c6fa4a29c0a9130c252532ab405fbda8e9027c094909",
      x"75e15dad637c47cdc342b40ec3836538a9f89dcf436a32edda134baeb0050748",
      x"c5733c733e9a788efeb17942cc805870c1012d71007924e08b0efd34d4e8cd92",
      x"4a3105f622e51c2ae5df0046fa2784b4c103a953705edbad73188b760039cb7d",
      x"4821f7d75397554dbbbdf1e4f3661f87cc3a8c742c5f0494fe488cec19a5f57d",
      x"8c358ed499bef9089a63d558efcfb4bf395bc51226705768e611db92aec2886f",
      x"f6f5f6140920dc6c275c0e49c999ec779b7861dcd25de17cc6a31ec1fc7c0c9e",
      x"5ca864d13e89728382ea3f1820018c8d490635c4a42ad37c790a8f1dde90b7f5",
      x"83fbefc06cb8bacf2904e68aae9b348b6c162f35994fca1f61a20455c985b920",
      x"5717e05b37211ccd02ea41917712b4eb9dc8aa454feb22d5781a0fc35046954d",
      x"2afd468c7add9f5072371bbdba113dde4288c3f27a2c1818c5751f2370b04a45",
      x"2e583d9eb74581c14983c7f4e8f5624e4eba9cb30a347b13179c472473f30541",
      x"4587c26d13f30f85e53b99a22b3879ad6f1661d93bace23419c88abe38710fe4",
      x"450da456a6e24e6aa869ead92add1f7519a9e966438ee903e7499ff19b90db4c",
      x"f140b15580b4509687e46007690c1245277563087004f3781c210161a4d9e6b9",
      x"2c41ab66ab933e1f58dc4f9c8eb664e4857face06f3dcfe03d656685342eca54",
      x"adf586580307b81705f8063a77463acbdfaa7b202059444e647184194a676d17",
      x"aec326b3e1722cbe37bfc2db6ac951dcafe66bc3ca019ee9e939a992943d8f75",
      x"7401d2ebc4fe9aec2ad8aa67f574c7f33b9c0a9bbd77aa7119df39036482a411",
      x"84d6f93384c9d419508ac82ef26182131e0f49ab90f49a3f8acec4194c8ee493",
      x"09aa78546b12fb0f2dca922b4b18cf3d5b28b3302e38832109caa341f3dea534",
      x"9453cef5a83ab81a94ba461b140ed86fd3653a52036cf8db412ae68dca82d769",
      x"03fac86748ed9f28f93a90daf8697b68fc3c9858672e542d8e1febb682422f04",
      x"c5daf1351f67601f714b3779b9703c9cd1ab85492e2a6c5089a67fec28089220",
      x"cda02b58f1a53a94d4c872481b574f36e7b23e62fd56768b5e5fa9fb90c0b1d3",
      x"67ff991c662ef8d8080d02b1b38190da366841f7bb7ba8d3a7ceeaf4d51811cf",
      x"db7dfd9ddf950153a5076da09cd901cc4539fe267092ed6c67a0947bae186d60",
      x"0d6c11dbd960e3a47d7825763aee6a8b9de8eaeebcda07b2cd766f4aec7c248f",
      x"ce900a06870a9cc1b39db259d016278d94e68f75a166d585cf463ad381bdad57",
      x"c8b63674d88c65fe6c12756a06b5147cd1021177e4eb3fc362f8c47ede1d6c7f",
      x"c055643bffe2479f7cacb9215b51368fa968474c22c451afb4abcf725652a45e",
      x"9ad927678e672004584cea27861c4041f95d8758b2de11a24fc155fc6af7a6c7",
      x"20f2fd653585d182c6bdd702a79d8546747832616d035898b33e51a29c3a464c",
      x"9737d2e32c276625289a6c4983153b3e69863887028ba63bf22f0e100ba82278",
      x"288d4e660feaebfb6510c516a1e377bc937e2a3f037c2e15f1aecbe0d7a5db23",
      x"cc55b16eb71227b7e22b00862915cfbe9c10511f671da68e6ca6b0f3d2a81f2c",
      x"b2916c891ac869c7af0970b28509de6d0a5df3fe6333246418af5a8e1817d7f0",
      x"9398d3f8cb19da1362877ac0038782abc6de6a69b8c600041b9dfed2861dbbac",
      x"e37f2ace0731a8bba73ad733fdd0b34a37c6e09242b1720ddeaa083bf565232d",
      x"fb9a79fa68aede759d117e32735bee56ecd1dcbc1fa55571f37159427c14b217",
      x"81e02e8c26164f986babda37e1a7943c517ede83ece6e01edef0706f7b5eebe4",
      x"7d095168084db925db4302eb8ef4d8252ccf2a87deb308448ce942b6cd629cbd",
      x"c17ccf56e0dc864f6418584c7a51701c83e3d7bcc8c83c542d1c375c99f4dfb5",
      x"75d9b5d3e4767e7f449932a5130381e160523786688ef78fe54f226e89fd2a90",
      x"ad79dded88d688f28376a2873fb6bf55c527d63ea99413ccfb7c3d0315dbdb71",
      x"3a935b846897a2ba3caadc37925e7a4a827c9a9383afa575deb979c7d0af3e6b",
      x"ceebb477e70259dd40642d1cd653acb259b89c85fdb53c2cd6878bd73dbf2dba",
      x"66df2820771b03fa369317e2057cc720678174cebc8d6e43752515dfaab21e3c",
      x"b9203e68b885d93ef954b8bcb8f22dfff78beb8c1256c9b446b0cac7523356f5",
      x"65e2f01712c6e9c41ef63ef7997445e0f1ca1c55e6ed287c2f378db0a3ce8c84",
      x"dd1e291cdc3e6664a7d9d82dbbd774f610666bdfeed7d0fe09660156d460beff",
      x"fd69a06788e59a95643302a7b27776521529346c898f0918e465721246978fcd",
      x"4b9a139a5b82949b385c9201152f44f8a0465343403f2dc91f06098706a2ddad",
      x"ac631893d2d92d370e73debedfbf5ff2e9723de2e7ac929258ee8435762e6054",
      x"ae896f9ed0a4fcf0d9b96d729782c65f9832a56526e0f2e0aa39db60e05f515c",
      x"79a75866cfa7371432401740fd8bc84b60ab7824c6fe490feb301ac956a7b879",
      x"d25800d014ed32b8e903ca686da46bf11220c0139bcab111bb519f3eb42be648",
      x"a34e2667c75238cda497994c3aa631891f5d027dc712fb9bee421415d630a334",
      x"de56708cdb30a673490f27d99ee5b72906b89c46fb305c927676bb858b572819",
      x"b735ba11d5df855aed152a7fab30ff59050b3516b51d771b018795e21687a7bf",
      x"f5a49e1c4f8f87791ba836befe4dcaf7c5fb5e4051523902115fe5d69625f53b",
      x"da481cc2f609134e3603b927d31c07f1e605a9e56e92accf3462d3a7c7f53614",
      x"d472d852fecfed51995a907efc9997e9d363c72bbe0119b506d375a9e860957d",
      x"8a29812dd56d90e08919c8a3f2bda9eeed7cfb7b402178498671454ce6971461",
      x"d2d2bbddd8795565c554d2f9c7679eb2f77628c5a8a3303777a0390ca3d9c0c6",
      x"7b21c04648f03ee05e3ebf28f0ae9f482128700e6d43e14540af57d36dac00de",
      x"9db8fe51f77310033dc218f2ccc0b8fb10ba1a6e662b707003b8c11ed9a2a7d2",
      x"769141152c83e06ed123ec2fba85cbcc6136cf3910c4d64f64e3bb94749a79c8",
      x"edb0eb980415b96acb1ee8f83bf30ed10b5592851fce549b38bceb7777e7ce68",
      x"dc86e2e3b9aecd7bb08b6b48e1bc436ba51ae9469e3fe5e233bd11bd8c8b2559",
      x"9be269f8fdaceae3e6c9d936d053bcb261ad15498d0aa62020fcaed3e573b3b0",
      x"dde5b7679dfcd1ad19a3d5c4b0852d71ee0360b79baf6dcfa4071b77d27c8846",
      x"ef0046f6a0a5ebf60ac7fe453366ea9bd11fce7ddf790711a1fa45170d61251c",
      x"f57abad5493e7ff780dfb57069e2336c30bd0f9a55a15c4bbb3b880195a457ef",
      x"7c267eb9348c5cb8dcb9b4c108b8ec77db7c93141938827e565f2ce1feb7d523",
      x"0d6521f6b93e966b776f5fe2a92884ab512c8a330868bea381535aa61fb09cbf",
      x"ef1d348a277c98ab4227d197c939c39be57ebaa9477ff0853f145da99885bab9",
      x"b9ac33c874b3bc6ea46a1228ac1dd5aff5bad77294a0a7a87f4b661bd9234c4b",
      x"12d5667b79b7764b4e90c59ba84ff83c1c8c92d6515c042e1ed05775de451f01",
      x"9aa88e897bcafdc71030363120b91dc7c779ddb31fc56b07ea0197eed4c2d125",
      x"46446be80ad47072ad589cce0965eeb4137052b9eaaea6809d2322b3ccaa277f",
      x"a83c8afff1e276266d24523c40c0442283bbf17edf957312eb4b5d0061322061",
      x"d0eb918cc6e38ef07860c19b1f8ea371fa2437349d268d9ee8af7ced6397a01e",
      x"eed3124a8a8830421b4ab1f6c3ca071983981076b6502ddf0abf593a939f9ace",
      x"10ee4693287c63ba8f915a7d7ef56a1875db6b641fb0f41d15fc215b4a0f6353",
      x"46d8e83e167a9214e87a2a5794942668b361ecb12f7e805f8097b32026d7c46b",
      x"9845fc5b5fa68f1b8969ab7c75ede62304c5b70cb32aee9c58db38ec862526d1",
      x"e7974fa7cf867022cf6bff3ce4c33747cb526f03ce01954f6eaaf0f48fdfcb95",
      x"bc81ec5402ae1628e439f1e1d2429c9fe8101c4035a8b3586cc81f3f4644124a",
      x"fe2802151ca55b1feb100155ec5e69db1af1743b08fa3a00e36f2fc9a0f996c6",
      x"288e5cd78833749c5c04d5500869fa76d33f516cdfcecf2496dff50450739d24",
      x"e353c23ca20a7e1d2bf9a03a4f66a139ad19bc842e2dc0c97d795b670674ef55",
      x"96059c87f4958053d70ddc4a647762b4d4cd76fcf7187b916b40970edf7b073f",
      x"9175e2b63e55a0030e3aacc81c0440e8669adc3c92ac5d4640157d4704707fbf",
      x"842c5a0ec925f8a106b4ed3c93dc5a8e30edf470eec488fffe3168e3bb26acec",
      x"420d562621070c82f026e74f8d3bc2feb6b0d35054fddb13bc5372c08a5e515f",
      x"c847be8e271d50c849b4f59674e92430cf90071746f583c3a1f6eeb06daabd14",
      x"85fcf58e0909784626332a5b2054e7c624bc447f74979d018b625982bd036821",
      x"8fde900025a569e4fde99576c6725a858f692dce39509e93535b491253be05d4",
      x"0eafd030122e72dd69a62c8dd76f0589f0ae5fb0d7c8f46715f9b38cb2c230a9",
      x"efe15bca85e50887c530e475b296d1bda4e12645d07c27f0b70230b2593b1697",
      x"4285cd1b8ab5456cba1afa468a27513245ed708f2d1aaacab5ebd48f9b755d42",
      x"2b6c80b12f53dfc9b2e23f5ed07dfe969e52b2ee5683ad504e64153dca1ead49",
      x"9f28abc2299c154553f1d3d18be36db12be061d48509567f2a78a29601e8985e",
      x"0e3ee857ebf036af8c3d1e55306cfade7cb46a8223f97e4279876d99674f51c2",
      x"81939db0d20521e796c199144d49cce366c0c300081b2b6df5110847f22f49f4",
      x"eec883be632751dff0b991ef1654cc79f10c0c8b9060a440d3cffc4a19ac1190",
      x"b53b716932f9e0ac0b3b582acb597d0b16947dff78aad3c8b62f7a4bbc4f688e",
      x"b8f0c024b56574365eda41e021fb7b5d7c81c18d4c06142fcec7bf5d5b66f893",
      x"eda7f29e7e40c5d201b4d3eb8543f0f9e03a32a1d9c8bae408c8e0d69c20f8d5",
      x"e07bb38d44ea2cc13532197a9140668f80063a46b9dae4a16865ab10a2320a23",
      x"5fe517ef488851b633b0348b8775087ed15efc91781b650e9b508cd76d887269",
      x"a0f45beaa625d01b61857943f2f38667119fe43e80cbf6e81050b9ce04f01beb",
      x"9bc7a921b7aece1eb4a6c194747ce8fca43dc0f51a0bffec55680c12f52b7cfb",
      x"f713ac0486533690dd5a1aa56152aafe879d56f6349a9fdda10cbd5624859e0f",
      x"916ae284118e0ffb8789dc40719549325926da97de0bcab0a688f333a214cd2f",
      x"fa86cbd17ec67398c01613a2ae669390b232d4d07cee15ff79d3e796b31dffcc",
      x"eb6df95cfc56231c76d16cbda6263c4148a3f164682088ee1e090c90e236d40c",
      x"960f67c8029d968fef756bbfc08927a03ede2fa118ede63bf5f43dee8a6ff5e3",
      x"4acb37eca34f80912fec911be41b9a78edda41c32603f9c87c6d7f61786cefa7",
      x"fdfc4aab3f4c1d19602b8394daf7fc3c8239e57faecd85ff065ade0841f28bab",
      x"9ea7791bc8f857284111b495ed7839ecf3320c79731769e39e833b68b82fc5e1",
      x"8a7869f943150dce6d7ede9da7db029e643a0913b7785f59fc1a9a9e5fb15f55",
      x"cfc57373734dcf40617c824b99d97a2f8dbba8cdf4a3ea2d57828f8a0fb2b625",
      x"d2ba341e219ae2e6db3b094daaafbdf09a38deb0cba33bf210e4a8a78e1cc120",
      x"43013266ed75cdc3ed69b541a50fcf6cd0f0cd2bfd3d63d5256de8099e964930",
      x"b57087f1f0bf5e5190d19c66a48c149aac0830531825cbc99947e7c1e39b6f73",
      x"0d7264458d0b833feae3159e0d858e193a995e35c48b7647e30dd62292284251",
      x"0c7384c51224155dce9b9ac20b1f3b3e2a3ebfd15e1cad77c2655bb74d8b920f",
      x"76218ee6b64f5dd35b463e894ab42742249d442d0102aff1810d265ba341584e",
      x"703e430b480ee011c28f50ae8f03d3e5eb769fb64a3505340b6209e2265a1c2b",
      x"d23d3b3c6a791af3bcf1a2b1ba003ab345881003174a6e150622e61d68bc564b",
      x"1e9439a7b76ebf782d4e3e0bcf17854ea8634ee5d55e69a6a07c9172b02e4d3c",
      x"766545412929fa49c8de8b86db7c27be9da0284d62653f7a6ac376558a5ba81b",
      x"4e59a0460b9569b2ab93c64217f78abae3b9c5e00e8fa4f33008aeec5a7864f9",
      x"83324dcca513afa04eb274ee219f0e461cf0a87c12a1b78181e70c9e3df79fee",
      x"6d3010587ec1d1888b67e2fcc3cbe8bf18db523b747fe885b18e58164300bd04",
      x"1e656b16b8f3c2b4878452b6a8276e645fd0c5fa97b5f036d220bee0263a740c",
      x"601363b54478e66030ee13fb9ffa16896d75f9d8c2d44d432b5e552162414caf",
      x"48d8cc2795092428155d5be0957c6660e0c17aaadf08c17a93d32d549eb03de1",
      x"264a5ac793224c2c23aa36257214f1750ca6b99d56b6586826bd935f01b23b47",
      x"93a7b7c8060b50009cc713519a728e66ff0d45ac5db61fc64a63b8ebfd0ab0d8",
      x"f89d1b5bfcce16bcd54d8438a2ab2c7405c8c767ac0f8c54d77972435fe097e2",
      x"c60499428d70164b6c58ad0faf483baef77d9acd1afff2f9763256b862fb6e6a",
      x"b09f9560f976caba5fb18df3c862253151875e57f33936325ae945175dcbe26b",
      x"bd816d9d420a3b183b5b0c4f520e9c66d3394b07ad4bcea49fe1d6480519e856",
      x"3369c99533cd53d44f974dccda41a847c4550769597760bcc4cdd1748aa88537",
      x"1f7c2e204761419fe845b0836d198dd81eeae5954bb1cb20c2175e84a6e6fbf8",
      x"3d1e48d8a41966dbfc2ff0172e209038155703846b7316b9e2e1084665abba3d",
      x"0bd196104b40385c31c524c2e7e9589846a6d9f55b610d6f4a73e6a5c3ddbcc8",
      x"85a05241c6280f7b81191344b15e33e378c9ef30f9797e2e3ad139d315a25eec",
      x"95ab4d303691188561d8a16619d05a8402ee2b7a73bacdc10bb2d7e2d7025348",
      x"0a758c22d8a86f1bd2eb7e440bcc236cf580dc190f20bb171a899775ddb1da2b",
      x"286c154e68bac72e35f7d2dd3f07090abc5c9d5b8c63203b41747095cd7ccdec",
      x"d8af9d27d36eaf5513a6e9bfccfd74133ceadb6a170e741fff15ec2994307da5",
      x"d7330dcb8b85866a9adbdec1685523ca96fcb79db7a29d9f3c14f00283a3220e",
      x"df26bd2e5cc09fd5b53d2e2310c18b0ddfc8c3bac3d72da32bf4d51643ba050f",
      x"52a331e7a962cccfe731d2cd6bb8f2e43ba8358cd0615456491bdf4ce1881ba3",
      x"2ca2b416c067d8a43a2e44750837310f8d49af08c6d37f8c00b690a3bdbb5219",
      x"78021a3583929855cc7801bc24596786ee5a5f2fa14c9b7a794dd0eebd76e365",
      x"1a74624cc387f9988b0f175f7313b5581f90fb78ef4d244347b19f3ca0d33de9",
      x"b651f22c8f04a38c493cb2746ccbe06960819c74cecdc1bacf63e1ea49877a18",
      x"ab18387f880637420f3f6ea8719a203ead91eadaf72f1c9002f892e53e6e5aff",
      x"a70e8e7a2775f708b04179382d0c07e738a5d6ad8d8db084b337bcd4e3e8257e",
      x"00f8a130ddb236adc942116173ffcc9ae8e0208c773248fe7dd0f0694cb1f10a",
      x"e7cb9d887c7de825e8df7c7c0e36bdadd3b966a03578b1cf90ae4abd40cacaf2",
      x"c2bd056b9b6b49304ddbaaec50597692d2fc52b4f7a237428d03530906b8a917",
      x"f8fc963f8e47af22f707dbfd3220ac6d36373fa857dc4b70bcb8bac226376f9d",
      x"42fa2a8a81804530ddb1141bd9e55992594bf637b84e4ede4e73e38d24654728",
      x"1d4d48c0ca3873b882d5b6017c853c2e0afde6a36a0c3674c621652acaabbc6b",
      x"274c3d81b598ebdc42e26fa387bd492cdbedab607fb3d90988da16dadde5b04e",
      x"ec303049cb59cc53051e19d8d9214ee843b401d0e28180cd18de3d0e5082978c",
      x"0ba02c34e87eba25a3336b14f20aaf9ccd80df0d38cb643d1e47e29b8483aea5",
      x"a8849c61a5b8867a5eaf1dbd8d5dc5f1e16199debbc07d5fea6b98e2c8e2118c",
      x"bff1a534ea5e9daaead92a9cdbbfd4671ce4ff2ed3aa1a9e3a8ae0cc21587b61",
      x"f53f56a5196d693724fe883fa4bd16d90e1728ef106a280a7f39162c4219e2eb",
      x"dbdd8c7d01be449000c2b76afba602c286676e821cd613ffd1e544ec14aacd54",
      x"4dfcec7160ce53d1545c4fc3582af136321030256af6904c0e99a56b59f3676c",
      x"8b8916b1212b1a6d95dec12e1b4894bbee3d64d7951d718f0ce20d7f36d689d1",
      x"f70287240621f7ff97210c8e57b5bd38334f8b67c3837f16b8dc95dbcd50ea34",
      x"932d891391e520ac689c674fd9b1c4f94bad00ee7bff4bd1ff103805e9156363",
      x"eb0ed893e5e79ebf1a7162f8b88668a14e51f1ac673d2c51bc7ca549136df127",
      x"5b6e5e4af1bd9522c99bc501db08e99e8e070f5f601eae75da7f080344940625",
      x"fe1255cf8daed3d79bdea79d94afe921f438d536610816daa38e359d190d1da6",
      x"043c7b4a10a763eed2d5d9687afe3cfc638ec1914438cc190f055215abcb091d",
      x"8ffdaab063f15fdd0fa3fc19518fb133bffeb5c66f9de60f7ffc6251abb67ef5",
      x"a747ccebd8c92f06101b2a0e1f8ab3de3df6f480351de66f0697e4de9d893f62",
      x"2a86b59e1409a6ad67fc774181a6c2a35799bceabe3818a87ba8c0efd6b86d68",
      x"7451f83f8b7ffa9e3cbe792cc0213e09d3b120e3b0ed98a8e730bf36dafe9c66",
      x"dab68cdde6f3d7f564689a3e1d7045b4f20d100415e4e635cd7e077db08167ee",
      x"fc48a8714e140582fb8ec04236d9f33c2718a4aa3a9dfb50670f520c4fabdb19",
      x"3a05be971b96e1dd01cc35efac1ab4924d9dcf3dfd24bfe64a6372dc519b282b",
      x"63521ea9bd0709d96d13b8a4089a9899556059daff075b77b5235454b70f5a6a",
      x"d3d14da8afac6cf374d407c6038b2a955325a3a32b3ca9c176c20b8b68718f04",
      x"e46c81f67c126734f752ed61c7c72ff8cfb3470de2d3217fff407c58b6f8b5f9",
      x"0432721850c66afc39ba6c08b527d510543841f58c3ff3b0f946c0d535d899af",
      x"e3fd40fb776dee1609a8a70e038f7727c5358129ac3874a02efaa50d8f85469f",
      x"00802bae51bb5aca389e37f184221b9085a7d9961b67eb9e9c3ceccfb6d4f573",
      x"9466dc0b23794b204834b82f72666227c05d889e0072cf35ffef161fbbf5265e",
      x"5f35a12b48e7ecc8ded9b51089707137599cde69a4561bca278ecfa150a64d54",
      x"f4ff48c329dfa927ac716426096bac284ad0d5d06ef13ec1607b74ec33bce8fa",
      x"8d76be94c09aa3a2492ad7ac9a8093894fb8174474759e69ae8e54e4e64b2c6a",
      x"fdae8373548e3a4f2f86118e731c8f8a1d72dd1c3e50e25b350909e20fd0cc1c",
      x"bdb4b9356c8e7fdc2a2cb228c1a38b56b9c7e772a9521af7aa36ca43b16ed2bd",
      x"086a72b7d8ffd0822a1802258355eb971b237b127a8d6f7a82fc493fea93be64",
      x"5ab37b4b940d09f701071fb3efadea0491c1a08fcf0979c6ff1f95c7f5481d84",
      x"23e494e43dea5da579dfae75ae7d01130d1418ddfdac574b7c0705cd3f358487",
      x"d41af7bda26ab146786cfeffc8c6c7a95aee27d6e65958abd2d3bf4d216beb00",
      x"7788d374dd9c29898f2a151e18a3e2f6fbf08918d2ed6fc5db1ee20d7326560f",
      x"a48b79069d87ebd4c90731894023c314bc341ebaffc95a87ae2b048a36270764",
      x"f73357ab07161f16edbafd02040ba11115860bad4d909cde5e1b1fc4cf7372d5"
    ),
    (
      x"73f90584c77fdd7138250a80efb8b3edd2d3dbc47baca054774b01af046b5043",
      x"0880b12f4a30d0618b40a3afbe51e37cdc0d11f16b66e3de18a4e9a0d235f534",
      x"a01574e0ae7fbc5a8ea6d6b979ef323b476cafcd0ece1c4ea79e250ba31da394",
      x"762dfb6898f2e3b6ae27271379bc0303c49880b39d1dc325178ee719d061a9bc",
      x"61999d76b91f66226305628a84b9b6535907e3c65b3b41ce485abb3e008277df",
      x"67f46b0ccc07ef4dc879cc46740a3dba82a105cb4cb97977bf44c67b5c33bfc1",
      x"99396dc62979d220cae60910b3845fb426b74763640d056e3524a238cbd19b06",
      x"5b969040f41cb7d4aed0dc2e8ea2346bb7d584e85e5529fb5acf58dd9ac8ed46",
      x"91bf14064bd361e88877e10607cb6ecd1023cde4ee0d555a50edbc80d7bb1bcf",
      x"767d7a2988da74d64ac6a66158c21f9114377dae343bfd9a6a7b5d10e1c26a20",
      x"debf165d11caad3d5daf461a4c50ef5c746c982ac54bd27135ade009b9dfa01e",
      x"bf96af5eb475a0d2fef8da6ed575e55070dc89a9ba8c2b42747895c9645ece23",
      x"9b520220ebc79c8838328f22626ed144d3b08ffbfe4ef39d6798d0bf9eb92bd5",
      x"1ba6afb677d8c57dca2006e16bf00733cb03137c30904de598062b9e4bf3a31e",
      x"d97515bb44700029519bbffe2c9a2bcd004bb3cb0f3e9c692fecb39af09865d0",
      x"1c91e7ccd034f29ce65ef3e25e818f482fb48a34118ea769cb35f06b4b9f4633",
      x"0548362758e92730ccc99ee4351f4b7bf36dc1b11264361db8c0761486a6594a",
      x"8b19d0b5e3cfe1287c5a9c03c1115c49a010697a7086baae630178aab44c9529",
      x"6fbe679379d1cc5773f615f08fd86554349af7608a006c1fb38e104eaff2971b",
      x"4b97ea36d6cb308c7b83266b8433d27a3e0c65c86e75d4af6f0841bcef2f58a0",
      x"d09a9c6be6c6644a4fc7350d4b1a73073623d5077288e9b3b97a7f19829ecebe",
      x"dee168c235da0a41835d35b5f9b68d82f98256c12c65d9498387ef39eefc04db",
      x"9e44de504c40fa33c0795f5272d9a3712a7fb834d92494e06a82718b685a02f2",
      x"1330529480ae75eb3757061a9df5b537501270761a154b309e3c208cf95e9ef1",
      x"b978692f889b61525c4f6613660dcf217202da21d967563fa524f30017a9b918",
      x"af8296d16138f1bc5e069425f867ca7a116d99beb8bc80936119f206f375b80a",
      x"7315c1b610ff0855b85f1e4b0031dee9a3e1cfe14fc852029b204c47cd6c341e",
      x"8d779c64cdf7079e2198dcb1d4ea58b1f76791dabe1e5fa0b741fc3178f0f3f0",
      x"2808b1fd06fe8d46152481081ad628e1d4b9f0ab33bafafb585777bf0a5dac90",
      x"fc84f29c6e3a1a060751dda57d27222ee6942ce47cfe62b0fe0d490cc57e823d",
      x"72eaa26e75c588007a3f18891450bebe7d18278035f8b48e11ae783bb1bad534",
      x"43f5a17ebd8012bd4ff31157733174d986394d1186fcfa2f21d3b140689e32d7",
      x"e339d0c2f7077fbff5471c1d1532ce68d7ecbe427829bf3cb70cc5ebfcf8aca7",
      x"959410fe1d7262d58b9165a2b18229d01894a6ca64af10aaffb74194d34cf35e",
      x"1885d38455fd0f563bffde5e5e60e28ad35e2308a656f5839327956b0d11b7da",
      x"286757f53e6177d403eb75280fe2fe17e9c4ee67a81115835414416d9cffb376",
      x"8b8dac9b1ce3b081eaf114d8270aef2d19fe6d819c68aeafd04df52fd0815689",
      x"c1da489acb10cd9f823b83e683c01f13f4d8a7ed069e824c1179daf026f8ba7e",
      x"6d25e9f90ef230caa403748bd112be3fec0396308b8a3ab93cdcc3464853f743",
      x"c0b93ed12063823e149f703074d2c1e8d5e4f3c3ed58379ff312fa3bf02093b2",
      x"21089a705353dfd4d3a38ba9f88a086e088174efb6ec18bb8dc14299910fb894",
      x"252b565968845512b205cdb3bd10adcb9c7a078f1c1e38000407b5f57b877e45",
      x"46caf1a2cfc7dca618b34905486c38a0d5f4bdef4fc00bac7f92bad5f682e1b4",
      x"788697146500217fde8bc1b3dd2b4fbb660efb47f08e1a0ce3f7141e2e0aa14b",
      x"86331e57a07d3bc9dc00d210cf4eb319f45fdb03ce4f54101ab12d718e034142",
      x"3b9df28779724a6c7d4aad0c265de6258c1362495e58cdd15aad419e03a220ad",
      x"ed36a0293da0fd762bea0817f8dd63f46d1e9e24a3cc9cbb40abf1c9cc9dc57c",
      x"5fb15a27d7419c033ac49a91eaf6018592f49437ad2fac55207f8a2e1417150f",
      x"6d24fb3e2fa2cb50cfd44d488006e2d25c4c8cf9993b960e9f6163c430fd05d5",
      x"406aea8153e829942b7b4da3adecd1208d7db92c04304451e42a48c8982a08a7",
      x"3c1a5d9616e552756733f5bc9981282ee1407ce0e644a2b8725b65879e5a20be",
      x"d7aace9192098dda72ce3369b39de40cd3d9487c22ffba9d650e51abddab20f9",
      x"2b8e76f15d5c7a34c31520decbb56a21f1eaf12499d757b6dfb26300ed773ee4",
      x"d7df3f73c6697f9449fc15ebe1745b2a8683370343e546e270783fe07c332c39",
      x"d609db00187f40a7b0fce31d6dbd1dbfe03592504a9d25633b64341241856b25",
      x"e1bbee27ee323dcd15f907ad606c96699dfa3967c9ae11b915d0321221ff0bf4",
      x"08ccbf319c6d57c0caf1fa59ea0525ebcc0dfc97a1356c0af350172a69569faa",
      x"c326c445b69ec342f8092b8c9a1d79856851a5cc103a99ff85c21fa4554cfa58",
      x"275e581a0e4ca9ef4f1f7d47751b842bb69379bc3d7031238337a0fdae543225",
      x"3b339a94aac8954cad7fc41972b1388e24a6609d71172bed15d6a3d09e657f66",
      x"49caf4ac6599db71b49a60cc579c5e1ca3a40a12161a0caaea151d1f067abd36",
      x"ee99b3c838e66be0847f3838f4aad09a4b7715c49973a9239a7a63d4f3cf76d7",
      x"1f07d647b2cbbe9c26297f6616888da90caa4e7a01bc53baf61f8eaf59871eb6",
      x"820853c985932b96b9df7acfc268c0843c30713c3953f8871a7645248ce25656",
      x"9f2a8fd734a68a0b4c057e5e40734708d4cf1f26cf3bb57561e39821958b3b1d",
      x"1296329c5061f36890dd38ca74c1b6c731ead35360ad4cf0ca3e0e319cd3c731",
      x"e9457b6146871c30123fbc3e69a7905299a3eaea784fa986674f411aaab92639",
      x"e2089901b1b34068d944efb07fa2e6796cf5ae6c8d66f610e8b551b2bd429594",
      x"99aa085173a1d01a1442fd0dec422332a6c57ac2cc6ca01e460a82471154607a",
      x"994c77bff81961d05be0b05c3a9e158fad58ca9359a879f02a1e89b321646873",
      x"401c7c2d1e974b3104fa53287a540846716a23f688b9fb8df21acdb7e7da21a4",
      x"587109178d4d6feb1936b4719c2ea4debe6a474cf7aeb7933aed8aff35dd7aa3",
      x"bda69b958fa5e3bc42a1e7bef19ba2015fbe887df18caab4637b4083b0850e3a",
      x"fb05060092a902939203d3b7adcaa180caad572f56d363464d72edf00f475928",
      x"5885863b15825c6137088d95eeba045ea5e89432396df35c7955497d676791a8",
      x"33ef6f2a23f5fedaa0a3f28ead2c7014a549832c1ef9c76ee9fdd564e5d7791a",
      x"4b467b4bd3edaccbaec55dfa758eb8d43c460aa0b815f353bfc2678358118ca0",
      x"07308f2ac4d1239a673242d2c2ac28653fa2d392fc24244e495b6ca95804a524",
      x"cb443a48988f02a7c26c898078b0418b442315d6d79e20619f0cf0ee64d8a008",
      x"aa9ce424bda67903ed88aeba32e06ce21f93b059e0ce5d33ea5ea741ea309d75",
      x"54488a35e3f56061e79510f933767396c63e1248c711bbf42e2c33d0971bd7ad",
      x"95ff6c65a246ec87a8da2350bc9fe62c6cada4980eb1ebcad9710bf4148c8e46",
      x"f9bbcd0837a29326ab6cbf358dc081f49559836ef20cb8c33881612df74b11f7",
      x"2189b8e14387556096cf0a257c9681a8c8b544c19a24faf35fb09e65edce2866",
      x"9ae9ce5fe9fa1753c246c310d0c803d28c453c2eeeb8ad1019d9e145347c7cd4",
      x"4b17d073532ad7858589745b1748ffcd424dac4a7944b966dc19735e27910fcd",
      x"86616cd33fdd0cc343a0c0466578d9a8455e0343599c58bbc020bac3598b20a5",
      x"8c3878eacb843f0549c4638398cbbf663e1f2f36ece39de63f00dc93a855b073",
      x"00862bb51960b8c033ec514f930f2679aaf5323a522bda8cd804128ddc9b8458",
      x"cf34c34f12a82964ca2843ea53da4bece22ab15085139a9adb6c2145989bac1b",
      x"b723063ce8c9bc8c5cc4acea28259c9d2e5dfd0d4486765f1c0564bba5ae0d46",
      x"f1abcefddc1e325d23ad2d300bc6f7898aaeb68e89a20a1aa8d80fbdb5a3c4b6",
      x"589ebe6efb2bac63e255fdad4dffaf592e7d88d27588be919504f5fa52b00761",
      x"fdbbacbea2f1c4630098f609bbe5de0ab5255f46b8431d50f7a68847de45b5f2",
      x"1643bbda355a4ef6c13a191a0b04c0f1fd718dc48296287ea900257d24641118",
      x"eda9298468d2ec1a798592e44e9c4371676eb96da117504a360566509298e604",
      x"de34ec5747ee9f79d51ec7411230572a9ad906fe6081c8e26116519bbaea9e96",
      x"eee5e15e55e83a041966aa272c0fec354d1fd79d726c909ae3dada106e06c831",
      x"678eee96fc0cc03b62940d99389985f21cf9cd4c2b52cff2b90971125b879965",
      x"6174e5c503cc8f97d2a218954f523d292523e99617453af885120b4034c8455f",
      x"b484929ab84d0827c266ab9436609abd91a40b57c01cd662834cbd84df61bd41",
      x"42177a417c8236569d6dbb431f48b979d73f2a086ca4ce0a932f695d008ea0b7",
      x"05bb3ce56f78cca569489c3d9959afe273567921ac183205d1a613ae50a684fc",
      x"26464a66091f92a481724c066e5e54e86a89da64aa88c9af8e7e664fecad4698",
      x"316ac3f38880935bbe09975ce3fe55268bd1ec24dd6abca4144d78942d6950d0",
      x"11a6b85b79af8424a457fc1be3a1ac3cb764099280c61d719fea9d2cb5fc2c56",
      x"a2ec39ec63ab1a75e8eb236f2e756ce4c684f35446834262d73bcceaa966cc0e",
      x"a714cf79bc6db7694975ba09636a9535ad8678c20db6f6f891b63cf61b6edb36",
      x"3c9e6aa790593c7bf0737250cb3f9a289bc87520441ad6b3fb089d037d0d98a1",
      x"d832caf820a8858252909924478f4c453bdb298d4eb58e457de0599cce055bdb",
      x"37eef7568268490e16ea57bdc1f6c4e59b3ff54ea4384bee54b2e19bd1d3a88b",
      x"3e2eedb5868e501f02da382099f087279ae0e7200cd0a38d4101d1111afac5f4",
      x"74aa78d7e2aeda0c0046333a76ee6fd47d35cd48da1549f7be82c47127e24ba0",
      x"170b394dd674f24375c8d3833881918852d20dfe99605585bb67d32450b887c4",
      x"89d788196e83c13d220216b8e870893d8a6e1b5c2e771f91384108982a88dd12",
      x"4050eea588cbedb8271b17627bd0c969a4a1feaa60a96bb39038054d6eac2553",
      x"c1044c520d856894602af6979bfcf609954fabd41140cb544a8247c9927d6e4f",
      x"8de5505a5a22a83b428528804340b101da2cda7198d2680029ccaee1b29206e5",
      x"c6d70047059833922c11461f8e07a2d1de4adc475296799366b94365fea3bad3",
      x"f90e306c1f5e265da34a80f4b1783135840e4511320ab557fdf12961c3dd6e9f",
      x"0b1141090e5dc8b3769e1024791e263ec7950ad2fae6ebcaaa232614e6f79c47",
      x"b2da6bf7b27c7931494828f1f4b2a345de51e5f1f6e0e92b4811a02febd81b0c",
      x"253d19b213de25c3a3011b0014b2f2fe55a160c8e80c7028427f0b623126b46b",
      x"2bb971f871ef5f9b0d9992eef1a359f544aaeeb40ffb9fbb94dae24ac304756b",
      x"0093807cfa31a5c5c2ce50805bc11eb1c3dc23cf0fcb1313c95f40bdfb63c3bb",
      x"a34f98de603008864d58230feb6db3d4de3a0f943fb217553e816c437bd8b688",
      x"b36e3fcb06efc79fbac1a030d78a25e9493dd5526e4ae5a8001792e6b4b68e93",
      x"9f59868026acac999e389602222b0180c6ea329983a403214d2ac58b28c6bee7",
      x"7ec41d864b92394bb6b6c13f7fd1874fc332b68e2d617c74aaf003f93bfadc8f",
      x"7fb9e8397e9a5d85473193fe5f07561c6109b78e1d5258c68bf23ea407339fcb",
      x"464776075eececb87cbbb2b1725fc49704f6bd285a08ce18fb6a40a3ee29ceda",
      x"2ac5321d0be7934c102b01a6b2e335f891644672b1576ae768c30d7baad2f63e",
      x"053609bfb7d64145f2adf90b7373dde7c186f6e55fdf9ed37a80ed5a806aaed1",
      x"b6b70b3d3b7b922cc28e430174b554c7ffa113892bc76cf0c491604a533eab0f",
      x"58190458bd041c31de3287423eeb430042b4cdb68879f0b360f5bb97a91dae0a",
      x"d12ad8f943ef7b70e0be2707c441482b3a67220c454041c22513b7ef898bdd11",
      x"169b87af058b9aad05ed949180b222f7aee61333e25666ebd43575118f74eeb5",
      x"7158e77266fe2add9b334c1526b092ef1775540898c1ac00e39ae52b9dab6e67",
      x"bd80f523f97372e3b41751d79feb5d84f5b389dcdcbdd71b4a6568437399c305",
      x"10ac573dd5017c3ad2b55adcc3ce1e3798128cfb2a239547c1837463181a9715",
      x"37fef68d599f9dc915b5f4ee2db2a1effd32df9b028485f73a66fba2695468f0",
      x"24a120cc2fa6181f431289387b892e06e060dffa1163858dd963082b21d9fafa",
      x"8751da4e0c3ef806ce2e47a73708671cc37856f3407365ba53fbdb96d410a185",
      x"e1b3874cc48eb5e92598a85922e76d20a1fa63cdb00c4a68d23cd0e1a80bfaa0",
      x"bde481618730de5a3a621f11d3300c96c41b8067377ba7efbcc944149b7fd251",
      x"7a521286f115370cc3d014ec87f2b944a0d1fd404547719fe8865a9705bcb916",
      x"3bceee49b5faa4fcbffd38c6fee36b18664fab38ca4a2962484e137224aeaae7",
      x"238655c247e32aa63dd1c3d5678d684983a99a7abcaad853695f531162da7888",
      x"e7906c3544b962f3d86b5a60b07cc445ef871fddcbe8fa0b0e9bd5dfd579c3a1",
      x"37961d0afdce5656f16c91e71bc23261a44f9186c14c7df967055c13adf4e244",
      x"7f8ccfd23fc341e235f6355b4e6aa09195d5db09768eb648b2a450c3a1904dd1",
      x"cdd645546998ca93574e3c1957daec2a849ec6658022ce2c2c02f93654cb3186",
      x"6fa7d489a62e84fd95be5dcc6836874b841cff408d6fbda237fe1cb6f82eac56",
      x"7a6069124926f1cf1aa9570ec36d3a401351026823c4d946ecae3a53e7429d2a",
      x"6796398948b26701d821f300e3f03e68659fb2d5f1b98f1e7c75b4aa665c1df3",
      x"758af2f1659f8529624ce598e7a4994aa9f5f7d2aca329c5e6115ea0dd1c1a54",
      x"0792fe19ac0f43fda087d8fd466f0b2ee84c07f1a5a2ef2ee05decfb318abe7d",
      x"fa49476418b853f42d9c564d316f7503fdef1e7042fea149a7a83c0e7db93e49",
      x"1d4f7cfed17e87d58f121eaaee3585bac47cc23cc16068f8d10f5e4354a35d73",
      x"8a2dd685dfed06946505340be51a7b73f6dfbb610b3bb480abca6dfcbd931206",
      x"12251cf55d31d6e2032758603ebe37f14f3255be64a2c751b3e85d3a191c28f4",
      x"c5e3fa325ad3637b110e3bbed3ac7d0770442a9caab5c495747f6933a55cdb89",
      x"a3b0c1e996a8a25b142c61ae04fb83b9f280c5a7087fb6805e972409ad29dfe3",
      x"32c00f1dd9fb44e668f8f61bcef07c7e1e15382fe92e0370a3264c8b2967de64",
      x"bfe14272840e11d0d72367d0e074607706164e7a2223afef9c208bf569d806ee",
      x"ed9934bba5ae91fee0a9ed6a381f37189c952ab9c15dc6bf13ddb555517aca77",
      x"9a2ca7f3ebb40c5d2c6d3911fa1f010ef6578d90173e6d19da57cd9df44bfccb",
      x"597d09ae2c6d98bf7990824a3aa369325c79f95feed8ac138276a7a5fca0c172",
      x"13d55fce548f825a6696f52fef8cabfaace78ef00a6854cbfd0dd95bdc1a4506",
      x"aa7acc977e67b9ee3e3e43b472daa89cd78a42fd09276f65f3b6adf014af875a",
      x"d8cc39608955d40bfaffd4933060b75a0e9b846778d1429df00b671b193140f4",
      x"567fa60c9ae9ec75aeddb7876f5aca8a348adbeb7d1d6cf48addac6acd389b7b",
      x"92736c36074ac42e6802ffef88c521badd2aa1eed73fd2b6ebeeed604e009be9",
      x"9dbd3882742dca2e93cac479bce879c8901666d32092de2a1684ed6b0cd80a4c",
      x"01e5580556ce321d90e1d9affd092bc200682c69faa367e3d26fbe26a3ef3761",
      x"9ce6f1b801dc78e277e4c172e46b109f1a08c4c26fb84d1692e205a2c9b2404b",
      x"d8ed16c0b3b6f0e3ee41dca2a9097ea59b71a1a75055235a7a2a8ff098e7f89d",
      x"cacbd4d13fc06cb1e6f891c9f1e84674ffd44c7326def61ac90cfacb76c0b34a",
      x"e8b0f1973fd0a7c5a8d76aab6d026529297c270bab54f1be4de761d4c9149a5c",
      x"3841d937471b8d9f3d1dd151ed35356e2eddf018a55d739f63e25ef93eefe114",
      x"bfcb3eb98f118dbaa9e7da0470e5b572276350913ef93d9914006a70ae89c70b",
      x"03d41c306892b8a42a29e81bce5ed9b3fdb344441bbfaeab0049b27b5b51b6e7",
      x"e41fc38087223c740859ebaacc385b9c6da789f71619a4cb05186941a4cfd999",
      x"bce6957661e6c06dbddb09c78920a247a94daa5127a44a98f8b35d590332bc7a",
      x"68d2831657f297e526f492e7f63823824fb180cbd9f7b879e5f5d54378dffc9b",
      x"0fa0e13594283c0015a0b7b4445026c76b37d87c68612f12ce38f649ac340664",
      x"5d4e11ce45169b222a30589c1590a1174adebb2235d0fef6dd39510a590a9cc3",
      x"8548913542649ed4e6abbab043ce22ca69a98298db0298ae878316388a678a44",
      x"fdfce1dc792056cfaf71df64e0d903c25d8198ef3a1aae6cc3778fa2bf778fae",
      x"8efb3c9d42c468c5bdc1ddab954a399c81db2b8eee9c4768f7ae3685d3b8fc5b",
      x"70ee5f08540483e36d3fab71f30b04bb18f724e04ddd4575ed9c6eafbf60629c",
      x"371e5521475b976b3a34a4c5b823f2358cd93eaa0a8ff1da9f773c76ba42f53c",
      x"ce780631a371fd6b3059119fae5ef2fc4cfca34dc1089c5bc2690dad8bdf7404",
      x"9143d93e6d686dfb9c980ff5acdd7cf33eb2e0338f1c5e3443e62647a6888af3",
      x"390736c10b315901fcf0f2e08ac9af3a93979704933ae5e5538a1af07d5ae20b",
      x"1fcc69e648922927f931def8f287eea377ec0fac58eb52ca2ed3693a13a5cbc8",
      x"71e8b6628dc78d1a9f72c0ba920cd84711cba9226a4748295fce1a5b5ad5e251",
      x"f016f80171204392b4dd38857f3e782e1eeb17141483457faf02ce28324e7217",
      x"7967d9143a5469d343a41937c32f28b1716a6d7b33ba9bb5716ac5b9914841c3",
      x"361445aca3522af94f804f3b5d88518f4dc30489afaec07a74cee1b490b2b44f",
      x"3600dc30d905c8d93cb35bc80614a34dda10673fefd7b01f7f6ce6e7dc180f62",
      x"cfc15e8e098f84e1179b85c6c403c95157b9164df835833f29fbfef758d8cafe",
      x"b277f5bfdc0a6eecae46c399b72360bde6589bdc0604dfe39f61afe560650ec1",
      x"12cfe40597d76669db5edb199cbe6b217d79dd6ca6f6727217641cf928229ed9",
      x"61eec12bf6b3b2c005d104aa615c79581c413d148eb35eca25e7ecef4d9724b4",
      x"01f71529b28546028d0ffdaedc9ce483a0075226a1793410108e93b614f7050a",
      x"bcd223223ebe54ee7ad68a80709ee3b614b99b42bcb9a7e871543d8d36eed335",
      x"ce9cad6b18629a990226b16a4699122f07578211407e18045403f577c0444bf3",
      x"79e0e3bb6023f34b5d5dfcdd41befd801ccf3d2d5653a39ca606bcc861ae7968",
      x"d3db3a55cfa6043c3b20946bba081c4754b670957be26d47e38cf579e9a01238",
      x"eefbfd973ecea26537d9774ee48ede678f3604b5d01d1323ad457f7451d07f2c",
      x"52b1a520419b52b62a4718f60104456ef1cea3b5ff7da2e8d1d5174b14fc1194",
      x"69214cf1771aefa9086fa9db8b7b36feca41678b912fb9340229fbb6f67f9af4",
      x"71d7183d80f7bc4a960413b63f04140b6c85017c1962d19a64d4409c8d8f7ee2",
      x"7c1f7eb6e463a5b3cc3045ff85a4aec0c2f3845628ec9e2f32202650fe15e3ae",
      x"d3db33a94f4aad49629c7fa950976c6bd22db0f49f079adf294d043b2188ddab",
      x"9af7c4f63c70357fb95b6321515f182c7d63fc68269ada102de476d60cabbdc3",
      x"4304125b4c5e061257dee85a504ccd79522175edd533ff83bbc35dc941a6ad6b",
      x"cffb3ed2ea2e1f98204e0fc9c1f59066659c3b67d560c4fda3d44953fc92d5d3",
      x"761d8d3c691044a6351f060f4fc2cc3ea23aa4707a5d1d1a0e7fc1c69588bc6b",
      x"9e4f1d1bf1173e067c6e657ab43d1a9144454c701d1a0b434d1b5716fd4e2245",
      x"4662eb0c12ff5932ca67f00f696a8b856aebbbb22096de879ad2fed6090ab1cf",
      x"d63f35fc0712b3db27f22b5c10517cd5bb152cccab96d6bf842bc24dda66c996",
      x"703f7921bad3147d6231263ee75e109cd5ce8866b8b43043500df50a38464e9f",
      x"133a20d320d61e6b400f2bbe5e0e55bd35407332aa244e762f5cb82c371cc585",
      x"256202bf528fbd679ad76b6a99c36fc03c11ac8dbb4e0154908483168cd26c61",
      x"c502457922216cf44abbb919930d4dc50ac1c26dd7760f618950040096a6597e",
      x"f71b2dc28ef7fe92d59e574f9c2efd761eb309426620a8bd876c0b0f43bd4dc7",
      x"ad85368e35b5b4f6c6eed8cdc3f0dcd5bad31c1f22fa2a6afef0792107169a0e",
      x"b0c31698987cccaf46b5090dfcf821a8371790e6df2f49eb1d0a7085e8545e05",
      x"7e9287060f204275bb4aa074e0d50f2cfd381078b160215e73c68dc03e71e809",
      x"d6f47a640ed3542f384a07cf60770c7c1dad54677bc3966f7f106a50c296464f",
      x"f4cb94ddb706b0ebd0d0cd6395b7d63ed4ea7a7defef2bb4f0238ebf286ed1c3",
      x"fd29b78cfa274d664ddb02fc81a382e9f43d871a944e186837e6f833149c0d83",
      x"e70195f5eade40087c6a984b4a7c155932b057722ff3d5513881454c99fa9206",
      x"bdd23cb16b9c14277716d061b19722270249eede962de43668663e95ce213fb4",
      x"6a65ef68dca6f09e2bb439222721236cc217c7f11dc17054159aa5d8c8f2e9e5",
      x"b0666c058bfb41e89b2da43c9e075730e3a43a72c98845232e675ab885ae8704",
      x"497a1b11cf670c3667d378c3803d3e777fa9352524b9017cf46dc3212cbd55c7",
      x"cc0091927aa74f3db88fa26f548cf54d7428a3f6c13c618f8d3f4b0c4dd53b7b",
      x"9740e2270a545159c406d11e106c19fdd37325726ae34818ac55e33232dff7a4",
      x"385505b1f00f782b05ddfb8c2787c13085f60ddfb6cc9feb0f55c9b4c87a266c",
      x"4358c2e0892a1ffc70ffa4d68ba2ea9c51f7c3643aa4fdf770def119668e7633",
      x"27f9d8d95f7777cf9459612e5b89689246902b67576b73f02d2c7df3d87a2f42",
      x"542aa6710ab4a676ba004dff2b4ca7fe2c85a5f05bb83b919df7ea7cf129bdb1",
      x"89f04e96399ec7bfa87d03b1147ffaf880cff029690a6fd7e254174ff209c891",
      x"6d4e7ce44c8e9a2718c3c7e88a19ae1e6724f65148a1b9158bc589fc20a2c7c5",
      x"e4e176f8d19ca19f68588494e8a7e89e6ec7bdf3eed00469d9f6b22de03184cc",
      x"3416175468a79928bb84218532c181212317c7a98d94cfd0f35abb345ff7cc39",
      x"7f5ce14aa4974db799c4dd787c135ac93e956862bccd52cce5041e424785139a",
      x"be0f0be596ba6fa9a7e6ddd4fd385d2a85db36b11ab32346e446ca4b60dfed9b",
      x"a5b4c815b522352a27964f6d7757c022ee8cd3b98b5097244c393640c6c23a38",
      x"07160123b632f345d4f37567b3dce74c6c390adc58cd0f4f3a9dfc6df9210cc7",
      x"0405ce3c168a8a4668c1e104ed05691458fe3e1d7cf9490e138ea01ef9f1c766",
      x"0a9ee9517483e4b55f9b9d666d626904b3c1fe14b1a3df9d63fb1408711ee498",
      x"1907135666feafd8579d458a4e9d617d70ceefc213ec880d29b7cd19af2c3499"
    ),
    (
      x"4744c094cc9550882e0c26b89c237bd0c20e20c3929e1ef4cb4369b64e430ae8",
      x"5cd7f4e1c7faf6505e3da96a95fd54dadc638b499aaf8d649c154c01345b588e",
      x"92f47a03b3e6ce5e7120a1402a61304aa4a92c791ca9a5d06daa3ced0318b0fe",
      x"5af1d338578bc4cf34d76b6f2ae28fc2070cbc6586aad59b4943c749bdd73ea8",
      x"c6c6c4a4635c5b573b708ca72d0c87e9e1b4c29f77c2cc75646b6891da900367",
      x"b5bba07e124cdca7a4f3d2a7987e39a37919bca46c36f4930e83b879d2a053c4",
      x"02bdf5c546bc965ce4d8813a6f42f4fe67ff01e518e6f16c1745e0f4f4af666f",
      x"3653a0ca4df25707f462074c9eb866c0deb09ac69272b7a869accd1ee6adff1b",
      x"092618a56d977bc2408daf81ae195e365c2a3b3a9021c8cebddc64b734dac04f",
      x"fcb16a60a888bda9aa7ced4f7199b52243011475ad571ca44ee07ce0464896d5",
      x"4d02c58987a7ddc7b326d2b208808ffe27ce589edc378f76402c22b2a6265381",
      x"1fa0c9004bdcb9fca9f8773d7fee8b10071ac40483a65dda3ebf57e17ef51ab8",
      x"db7a9f4661a32e08dea6a4d1dcaefde36022685acfaacabf84cf256123293d06",
      x"a46095bac0eea4d7cf5f510d19827a0673af4b5e96237b995fa956803135989b",
      x"3f5bf958104b9bbbb42edcada0b0feffa906665e543dee789f419e970d1def23",
      x"4fbef5b9e3e22940fe100482b5b13eaf8f3ce74314c7e9e84ff2f4a2a73d2941",
      x"38c98aa9db1ce86ddadd1bf413915fec3eac219bf268c830882f20a52e22799e",
      x"612889ee947990d7a71435d0d7c7f93c043cbb68119f0004149233b14762837f",
      x"ee8d0acbf0df6050313de33a8f4d67df84b00d4d5194f1002e5cf475d77bde54",
      x"f4e67b7bbdfe04198e377a768836c53981f7499b60400125f68e72f67bf2ad7a",
      x"cfe0021f499a3849dbeeae878e9afe7bfbf28fbec8475a6b3d618361b13eb17e",
      x"a2c809a958e23369d6d7e9558c7b463807547f8aa99d9acfd03a75aa8a686653",
      x"6c3b91c124dfd03117b4c1d7336130c4ab40214423ed0b731c65ce946b97577b",
      x"da3270e0c8c33f1eb72ea2442c261b774814033a6bf418aafeaeb7a625ca1e6e",
      x"e03ef6a12633f089c8026d799996984ed1117e42aec7418670cec867f56dc68e",
      x"beb60057aa1d1e5b2963dfe243682a56956cb969b94d3e41ab77264809b65f80",
      x"70107ceb92003c0993ae5198e9372cff992334e44d6f26418bff97c32957d2a1",
      x"53a7836b6a3b0de9d1785e43d43dd1dce7f6165bc6aca94bcef407a11e2b0c71",
      x"333ad7554c532a6ff6e03ab80ab93a516606de4e8bab00ca6382adf847cf96fa",
      x"686a64b3f61e143c676ebace077f47bce4b97e1828894023a07907a32635f569",
      x"f6be2e6dd11dff09002582bf7366c21d51f2f6923e8fa81aeb05b40499c2c167",
      x"1bd1fc082206d795fec4e2b4d3645971e8951dcf0aa1c030e1f12520e65a5cd2",
      x"3a741229f45554d2bc7ee2789ee3d773a6b2347c77a4fafb98d2d1efe0b8002c",
      x"81e52c1e027ddf5187454b583bcaf7748ca24a1c82c977d4c3e98afde982c9d3",
      x"762b8cb2b9840424af4d66095ae5ea4c026255dfc56c8d79fe32a6cb463fd8f0",
      x"f0206fc5ef048629741e3fd8f61b45c976cc2e8dbc8d265d2a55092c62c6563f",
      x"5f46d5a6148adadb3d89b1f821ac80336ca2520c3cb30d8f1d72ea8c40ee3869",
      x"2875b8f70f1435f35f616d15546259105ca7c3d9b1f1cb0fe260bb15e05508fd",
      x"83a252a9148edcbdee7ed2752590389f065a1d9840b29d7c6d1d5758b54a6e88",
      x"59923b16987f3f96775010eaa84ea8820920a707d53d59b1e309c0677154caab",
      x"b0ef28714b72bb09b893c989bb1213fe4474d18d04210f80459da0212883dda0",
      x"62e574c953e057273af206c809f8022612648b96de721f957f08bac60a74902c",
      x"acc7c3fbf079d002d97a14032b3da7da7e9f2e612bf68687daa582ec902e2811",
      x"f433f10e10e3c0f91d377ecdf5d8ed0a0f13c59ad5471acf3e444bc68a94dcb6",
      x"737f95f69543fc8d02452ad13d77a03b0b11c39481968651223c65826adbf059",
      x"38d3f5f8798ddc1d3b6f0d48d1107a017789302e81f5391045b7d3e4e3f9f7f9",
      x"b44285e1074ee2bd37cf73d0096675a33975ec47d08ca413c649e3ff933917f2",
      x"269030facb35a035439051a6a6d13da358be90c7e33312d3bc5053a6f28c2c5d",
      x"805ef66214e5a29f350af86e8f8cf0909e072d75b745ce674b197eae5ba6f8dc",
      x"a24b91d4306ff71a4b0963c72d83f0c1bfcfc056a96d5bb55851ff4a982769e6",
      x"25814e74a97c8ac6b7474d95562b4c16cf3753ac1649840889b1371a14f58fff",
      x"d9c489a997d10ea20189ee7ec96d40cc78a60c379132dd24982eaefb41889749",
      x"041c8a212e811814bd99bf8a28e35ba2dc437775f0cf4c7f99040a9183341e0a",
      x"e23333d636573d96d378bb1ae775e30b84b24eb1524dc1d5feaae2f73bb92fcc",
      x"7f1faa6fc08a16b09c3daa923580e4d30312a84139e37bbb30965cbce73e1d36",
      x"fcd5973e50d52f69ed772192ec12def3bea3e6f4c8a1c1727b8f3fad3af11d26",
      x"275dd70a4a0c0313f7c9a22cd76f04a48d536173978769ae369b878786c3a363",
      x"cd4cd1e90d8f5d58e1ac4156644f78ea7131ee28469d169dcf9089f8e1d3ef2b",
      x"1c2b80ace817e40d44198b4881d787517066fd992940a3765172ac9c6351a276",
      x"30406d656ac0cb33a1a457bfc22cbb6c84d3f80433f8613008e24e3266098460",
      x"02d045e4069b8e801d006ac51d281b97a3e153a6f9b5e3019531814854e26c37",
      x"eea1b56f57e14f7cdbcb3fd2215ca7fdfdc577f12f04ba574ab5d4e1b91e1708",
      x"b5603425d557e83a3bf25ddb84022d75bf8b9b21fbc902ed3c0f900c01c5efec",
      x"b81060ea5005abbe3e2451f59f4fa1e345ff6471f7095f15d1fed4208a11587e",
      x"736bd46b62523bf38588092636df54be6d1fc60bd5add6ee88f1b80be74d3b94",
      x"5d37838067bfb87147172cbe9f958c9a0fed42c7e8b74ea4a35332b1ed586861",
      x"794165ce497e3f87b472907e61d1d1119863a287a3b6bceb7570a7e816189815",
      x"46838e0711362812c1b11c9209ccc3dd49862456bad196a54b8ff32617a2de41",
      x"16f62b7d9fd03ab70512ad607ecf7af3205501c7b75552888cef2aa1d96d136f",
      x"1e2115472d40200392b5269c8adbc2a28aba53a5a080d9db13c34c38655a4ea9",
      x"76cbdc3d9c5cea7ed24616fdf019975d95c7a0eb53caf9a9b5e38d855cfa1b0a",
      x"21187a5f0b0f4149e7d2eb6812a63715d6ce249da693ed776b1b749a7a8a3dc3",
      x"4d22a90918c29df96752d28205e7f39192af87f303194b9f069edcf573cefaba",
      x"d70d2e2b5af778e9c7db5e0ec6318d027701da7059871081645d39a42a45fc45",
      x"337d2ef77bdd3b272c78fb1c8f102151f0e5545ba9ea9a62e0a608625f70c34a",
      x"6712a5adc83242ce31340815236328444297f0798c16b720df26f3802d8dffe8",
      x"8a8e8a19f4e90629215fa453a6c523ae60fca3b1b4df5e4d8b7e96b219747f42",
      x"e6e4b973498c28880af814cc8c6480fe02ddd6d150fa2d6d96085e6421a7bbc6",
      x"2662ef6d66f3a3ace618c1600f45c74b223e41c9bf24fe162fc14210e7ef27cc",
      x"06de3b2c6469c12248debdcfb04987c97414035f5bac6f71d69f6a8d0bc81541",
      x"882cc08c91046c63f9eae81099b3a05532c4a588793ab283d2915e81fc900f30",
      x"aa4c817898909c9304852dc6712206abc5d372fbf227d957c82610c50cbde2a6",
      x"fee2a96aa67d842068201843229292cec8f6a0864c91ac595d888f55febb8bef",
      x"c260ca6f72d4d7c41b251a98d66fa06c0ec0890bd9fe88df4de163ccc043bfd1",
      x"e023367497e33bdb795e837aaaed5f63e2053cca56d1ec28b8f3e4917f1dc7b2",
      x"f088b1a2ee6a8736ffd271745dfcf3e1361f3112826e0db8377307c2c730afde",
      x"20c7b73c5bff249c1f1b73250720d1c3e05eae99c45da7d484724cfb7241dd2f",
      x"3d2e7d5aa600f9ecdf255d50e4aebb11be57511caf4ef94c78f20c005ba4e9bf",
      x"2511d8be84603cba63d295eea6d351f639775306f45e26c266ff4e09c8b11b9e",
      x"4162502bb6932e7136c052e919fcc2ad1167294eba783a4daebd1e0e2f12bda9",
      x"8c2da88b24393668182508d4e48385d62d3d0e8c167bd13aba6ffb91d62a54ac",
      x"991baf6a9a1d66e34487c936decee668735287e2c2d0b9687f1fb637c87152ef",
      x"3eb733e150249cd52f08d069329f44f94a8bc6546497e05086de337b5b8e4f18",
      x"07f13f097bf938ed904d006929e2dd7d1d9e04dccf479e6479cef1e64ed851b1",
      x"0a9ab10f21f7e92cf1b5bdac4322f405e804840eb7cec0f8807f5b42092d4e78",
      x"b263d6542da0df8248ef557d9f0c5b669cca1c69c0cdf96ab741ef8ef3e7d206",
      x"ee188cf3bdca68b5ea2ceff5d9b918b97805a7e172241db2c44bb2f346a70678",
      x"626f958a2194ce3ef446fb5750c6ae9de30a5ba6d5310c11f3a5dcb2dfe70905",
      x"280b9377062d951feede6352844c96cd511333f3252810eecdbc9300ba676c7d",
      x"93f29ccd8875bd424ab8bca69a8d247b1e52fe551b19a77ddb95a66c504f0984",
      x"7aa7b45dd5760ae93d0735d41d1595b1ab49b15bedd34c082f6fbc7007aa15a0",
      x"413cf54941e08b35c81edb1a1db7f763288efee6dc3f6d03260eba2159f9ff50",
      x"05caa658bd5df974b4b9bf3bbd07423fda002130e6a664d6364bb0d94112ea42",
      x"8feb3ec94af254aaebd5046be327e58e75b326b5a3bca5abb011d6531c9db83d",
      x"067f1c7e53d49f406d23772d04c4dea0f6e6250c7bcbe8700a104bde3f34012d",
      x"4fe6aac632ae4599524cf264e6f36c407b52cc50a261ce4462c9c789a825af18",
      x"4f2dd419941a8ce8787b8328b39b22d116cefca2d7dce8685596bd66055e3b4d",
      x"80c6560f13be737068e671ef3b706ebe3036e1458fba7a356d09dcc280696aaa",
      x"44d4a682a42d406439951763651dd5c5e7c89dba2ff5d9891df5c8d9e4fcb636",
      x"0d78974443e4b0c758917114d9949f5bf148c6b1cf035eb4e856a3b150069a21",
      x"4fe8912c69b88beca7561164dcca5f5cff1bbff3bf17ad0b1cbcb277debc0013",
      x"5890e761d5ce6142b100a848ff5e4e4fcd1cb95cad743e90fbd20432dd71f181",
      x"95b5ada0c0a0b31f8434abc093be303785b921c63bcb21aa6692d1187ec4a1b0",
      x"d434b50934e004c5535c85eb111e5d1bce9b0706bb54ef1b96d2b1bc4ed9ed81",
      x"860d3347be5367a66fa9906b8f8f39b22390ed1eb4e16237e03ba1e1126383a0",
      x"5dbb8f5d7fedac9da84b7831b73048b4cb3f768aeba08100015e740312beab17",
      x"19a6f8556101734432dbcb46301c1dd9d9ff9ccb84086946cf6037727ea35e11",
      x"9896f4159aa7ba6ccaf6ea8d11b3c0e9ac8b05d56fb9c970a27a45fe90104f5f",
      x"bb6e78dae9b3af51c555e4b1ed2b07f5fb03c7af14fdff9ac6d0bc62f7fb2947",
      x"03da480f27263cf67c80aafd8666bcbdc55a4613ae02c0127f4498af4640d327",
      x"cfcb9703a4d312f88fe7d11222c4890535d76406131169cf56fbbdc1ba619491",
      x"ba76a47a504835ee1e8727e2e5fe3fd4a738449565e9767eb1d9045bceb2c868",
      x"4c50e99ec2a57292a374dfa1171aa107e7404423f6d9d6580a2a1e967f4d73b6",
      x"e43e392a84d031e13c7146e2b2b8f21df172f051e8202859a9195b5e260a772d",
      x"d4a20186f3fd4b51a76ae1226098b256ededa213e09e740223e561241be86f98",
      x"147e55c45bce2033fc3a3156e547b31bd47fd52dd0ae99285200cba102bec833",
      x"dab3ebcb2a9de566c17324a9d654e0de45c5eb582d8bad90e4626059bdbd228b",
      x"b490256da92183465032eaa3bbe77b46dda339581ecb980e0babfa650a4c90a9",
      x"7cd9feba22bad8b58f2f3e8eeef6436b36198c6368bf37c0e72a81ecfcf72a7b",
      x"b2785a2864be85aeaf63455492e7776c32b79892ba722f0a397ef8abf3a60591",
      x"55711fd0667b397ad5a9865a227c6054e4ba3c05d297c6a9abb6bbd364719c31",
      x"740f69650611bd1e2b83618a02df502545e2754586de51fd43e4a713c78d4fd6",
      x"f40312de4010fcea19b57f44068b6601fefc08c88d88bd8e40771286a600f9f6",
      x"4073c2b600720bb1ea67d149d367fee7b45212ed392eb78fa826df791d248e97",
      x"61ea17b25ab582e1305fb8563472ebef7d5d22af81675578d15ed05819dc223f",
      x"2a98b8d56f47320868d2081236a79e938ce77f93f535293bdc3c1b39dd5dd55f",
      x"5dffcde062bcd17b1cc79ec5599a165fe022a35e7463c53e05848b2b4c80849a",
      x"58b8655bc4d1b3a0ebba2987de27b8d843ac1cc635519524e20f9a5111a43e3e",
      x"205798f40dc742d9d31fc21ca2ea8c760ae2b5be3b474d8d7ae3bcc8a674edbb",
      x"1e33f56daa9bf981d971b77f50294815ad5170936a30b82083f2570445d51c09",
      x"49f373f387634a3bb6e40d74e1ad456b601fbf963e1ec2a11d7854b3f769e30e",
      x"610a88a966c56780280a3e347c49bbb7a7b4dc52c0cf684c90edd6cd306f5fc4",
      x"cbb36e26303f3119238de50f9888585295edfe6916dbeec8b18de7b8c734f0f4",
      x"fec5e95e356b90e8e65256df7fcb7e2d0ffa99535a806868f8e9003d48591e16",
      x"0313ae3a044baa38472a6fca7d1fbeb09b95abbfd764fbd710048cd6820b6333",
      x"32642e3b953ca3c1281ef88dc68d96eb8361be18797a1421167a37455ec0056e",
      x"36a731af0e6482991deec347e0b4cdfdbb148eb52c47fdfa637fe3f525e33224",
      x"d3bf06470cd2ebb6e98156396da68a2377f6b3aa757ff73f57fd0a1633593383",
      x"3ae00cbb6a246592025b5a3a5b2fa2746c1633578185f17b694cb337d445251f",
      x"f5045040ff01377a9b7690f48f398e60eb5d5847487e4dd9fad6b129e4cb2281",
      x"825681816d0e48b49e769a5304dacfbdc928aa1947ee571157408841885448f7",
      x"9d84839e21ac32dbdee1fb900ef23b417ed947b49725dbf1324b156e4697f8e4",
      x"aed9ff30798b9f03aeea2afaaf765cd2bf25ba25c28e142bd9cdabddf4fd57fe",
      x"3ecee88e04abf341cc42a543297a126c7f98109bf4399d8ecfc5a4f97de378a7",
      x"087b2d37fd547bc71edb4afa3d16ba7cacb2d9c9974cfed3b259a2a300336904",
      x"dbd7ad02657ca019487384f84123462aa2b5726aa093054388633cd7e8b7f102",
      x"def5f839bc4ca7e229dafaf51884dac2101b9040a3ecefadc87f3e786cc8c2d5",
      x"b9a6f09cfbd35296a7f6415c5fd24af4a9471973444d58acabaf9e7740170138",
      x"0c6207279c2fc5a1685ab8b88c9148a1abeacf6a7a75f86e601fe2bd14c9c356",
      x"14ac84a5b1bb635cad8551703b83ac8974884279e0fb217d2ea1f922f078a6d5",
      x"275458b1f57704a63ccf162ac8d1b96b61b3f06c8110b5a7caad484d82994b42",
      x"c46ca1fb0172d5530bc056c75b52924e9f0f1819a45db2a2d99ad772cb90fbf2",
      x"433ad43134fefa92fc3c2b1d9c7199a6479c111dc221427e5845dcf907e3eca4",
      x"2ae7d3d8df1b97697a455d7ffb56c59ab9f58585831353c89c210e830461494a",
      x"f347e8c9c82352ee13a113b51a1ca64bb839ccb61a0af1b0c5cc7c7bd34a1bf3",
      x"aa4a2f50796f514d3c3dd2b1a42e3262001d37dc2469324fe1d32ca030b67d9d",
      x"40c1def9da2666e38a2907706e44ee76930e08921ed1f8a2c37069c1a5a8c69a",
      x"cf513643b16550b29693072058815822f34f8402e2ad8ac6109b404f5be51f9a",
      x"4209d0e257a8260dbe417d3f0927f2f8917921ff9c23b9d6e3c6d8b659658cd0",
      x"71ee3b2b1be51d1ac3e28da49f3ed8e634a26af5fe6992581939510df69292ba",
      x"37beada39464dd976bed8bdb2b176d7fed7d81427222e9b325490a7c63115798",
      x"10f8b6727887dd8b47cd827277ebb0566ccbf134031ce28f5ab4ad700a1d5784",
      x"90cd65b5ba5ced9c5f1acc338f342f42d4ecfb3709e68422900c2b77ab6ba48a",
      x"c308ff25bc90966ba815526b49b6a0b2e0076e39c693965eb56e45bf9f7842e5",
      x"99cdda00d23d14fed14ee76b019f933585888a0c9de16c11d7292b6923216530",
      x"060e390b4f2b6af0b16461c969f6754ba8d03f5642949f25ca1489b6185e3ef8",
      x"70068f7c283d4a09f3d168bba763a4318e787fb9466051a372c1914a259f37e6",
      x"758d6fbdd95c4a68c86f74a8a59abed6e680c6f2234ee91a69eb7b3d27a6c164",
      x"f8f6476dee4d83a26d05c746c5c07bf032fc1532198e9b6d26938e65f4bab6b1",
      x"cb7ac64b10a72d72e7a5dca7bf8c420fdd5a5a859df7ae955de28ca11e26a18c",
      x"e3115c57407da44154abdfb51b14d567bc8e4c41b15ea69e016fbc123a95b9ac",
      x"7b4c89f252ad5ae3f3b1467d4498d014d27923b0554efaadfa89cc19a0a7b0fd",
      x"f97f52a79d09a37b85c434353df6751623f648271b0be696f343c75502706443",
      x"14453233ef7d42337d76c98d0edebed57bbbb42ab1eab50287c7a97da5bf74e7",
      x"51c53de6afea1533ce48fb63956d7efa6bb8e420f2bffd3017078a47ea828823",
      x"a05682024396d84fff3992c258fc6fbe5a1785197e480f24df995a26d33e1d92",
      x"c06f2e0fb49e5e26fd2ed6824e343bd849aafcc7c3a33493db73233140ec0b38",
      x"13d3583bb8538c61a4c3b1d4df5e1cfdeb2c11d3ece9ec354c1cef0f89a2538e",
      x"3ed18d189f230390d5e12b196d97b46ca0f36fd5bdfc95026d9a207741adc444",
      x"6cecbb90181b75d2a3ee0e2d6677d9d507ec8464eea6b2e13cd376f00c7fcbd7",
      x"ef81a19b44d8fbd3e0641e7f31f980e115690921a7151a2210691ed0ffb3ab06",
      x"cbd4cfc067eaaf815419e2d2627bbe342bbc1b9616184f5247caf499da37752b",
      x"4353ffe4a2b2816d13261877c02225e0e228a673191e39d5f58923d5576f487b",
      x"d722015921895b26c0556c7911927ae98d086a1fdca6f7f66373fbf4a2eae8d3",
      x"da7732d74350deec6b3801c7f620e7c946ec704b65f0bf7080caf3a87c001133",
      x"4fffbff460fa5dd97eb712ce7ca241f0c7d79b4d95ae443741a3fa69ba57adc5",
      x"88594270d7a5edad83c43a7e6537a8cb9ca67a41b8b970b75d692054d8679460",
      x"ee9a3330d989c794a41a2a21bb4c83376391c57b92310006364d88bd86f86715",
      x"7c56e6852db07a518464a1cf5e7c2ca7378de4c65525d2c49e53d56c5f93b712",
      x"0d13aec82c85ece0b6c3d8f8954c0050f595dff1ad09fc90a712575695ad4bcc",
      x"7643281bc79219ea14ccd1c86f6ce4ebb43a79fe3eed2e106396557ee60f9d04",
      x"b9e22c2480092a4ee9ee31beea3268e9f829a58105b4dd93172501f301c0ce0f",
      x"9c0929b5a413ac7090889709507ed5c458f1e91bf74084be8876e00e8fc60719",
      x"4d442df1dd4c30ee1f69eb9e52d2e079bf21b3878efc0a6131eae2fd199689f0",
      x"8aee4533307b668214590ee61bf75baf8a2d4f12c6ef1b72a733f79f9dcc4aab",
      x"b9597b09ae79e5a72bfab14354b6aea0b0653885cf293423e4fbd86ccc922c60",
      x"f6b755ab16d705cb0665d46f02523c30b7a41f19ec435cd7d2757fe74d2d02e6",
      x"3f96523cf849c9e58a8ac2bd1061008f414b71342e280bee9009f88e8e6b0e53",
      x"d5132aef70136418ba7c8931cbd695a1c35e2168ae2a42b7ea337d95b2793f35",
      x"fc08f0fafcd9aa3691def2cd5321ff40d1d738da527f2045c7ac374ed43ab2a3",
      x"47a1ec796f3520879dea592e4f47101fc857cba18135cf30d8116e6de846bde1",
      x"fbd73b0300b174fe381dd20930932b7eb7a30878edfc7101a3966b36fd9e4632",
      x"6da78955ab8e5efbef4fcfa2533d19ebb20a1684c7027f9e858f473e3eb7d27b",
      x"b86187effde8406ed5033b6a39f7a0e7cd533434fc5cc2232e25dbf27cc1b7a5",
      x"4895982ccff2c19e155104bc4639fdbe1b55390b133fb3712e1c9156ce0db88e",
      x"8fc9d38e80a12590fe7165bd072cafe26465db4ea0f827aec5f0533844516e5a",
      x"29bba16e083764d638889d53ba7d3c728a0bcaa19231019c8ea12db78b794044",
      x"0b8f4d8a37c45ab5ad4afdb94b135b2e0c75a73d4d6695d6f08aa45908e97ca3",
      x"7a27ad3aab5ddd6a1a5f431936ba4130669e2dacb85f6f38493446faf4b8b19b",
      x"6709d50e7d09ec8be63f637431a2ed028daa752a307eab6840b277d08bf57bfb",
      x"ce62d2eb2d0f065ea0b074583107ade7ea7a64a3210dd425c63eb0adc3ffacf3",
      x"5c7fa3a4360f1cbb91d3482f32ad081429bbb8ac6b322e8d0517af285011cbad",
      x"6fb3deb8d0a6a6651ab738dff1e59ef9d6641d397897ff53cf1a1aaddce3d538",
      x"d3c228f854d23c3f1ba669860bfe06ea30562336132e8765a8233e1705016cca",
      x"417578e1c40848fdbe2d42cf845255d2f375bf349ce5ce9ed9fa9ace21dc8cbd",
      x"83aa32628f9ce22023fd366ad7d1e11755e154bfd9e6fd52448dbb010e59a482",
      x"c651d6d59aaa7ed6e83ac3f9ebeae37236d43c97a4ee7ae555f6db9ca50ddfe6",
      x"352bdd5f785a5255c37da1bc772619d6700ac9b49c35856dc1bcc1b251ed2429",
      x"3048fa6d5712eaeb41d6e13d9c857640903d9d2c582beb14f420628314356794",
      x"eefe6a35eb23119e05795fd5e35ad484e3201a4591f5697967aabaa3584d1f1f",
      x"f6dede3c0334845fb583c7ef0c0111be08caabcbf1be65f2fe6946d6ba3cb653",
      x"71e3668392068579008c755f18356b4e20afe2827833a57bdb2132c84716a31d",
      x"465a9904e86c9d8432b8d0f2480c429eb5becb6d5e437d2553a2fe70796eda58",
      x"c545b67f6b30ccb9e94f68145a1cca52aa551ffecb4c1319806747be273aa128",
      x"d5bb54495691010cc64fa0a4c03e31888cdc73a9fbf535af8d4cb33735582a53",
      x"31778db08af296cb9b1c90afb2d7deda6f227d3715e7f0e76f96c55a1a5999e7",
      x"11e73011c2a6a6accee55b00e7bf4ad24f5f937775408d585a3271e788e2347c",
      x"373a34e8302680e023e4ce63fcdc638f18aa9c7b1061c14cb5fdd9a6b47634b1",
      x"f9d352bb7ea1badb4916d4b7b19e0f0ae5350997a246f4a4e72a36c9572a985d",
      x"f6122ac8fdfd4222d0d8a2f456ae5ad7e830f7b5130f2e48ebca2e771721878d",
      x"24f4b3e2a6a612a3577f2c69e89198be173c1c17c045889a6c4784d258a2575c",
      x"8014d0b970e27ebadfcf2e410c28757c19aa65927f30bf1296d43c8baf881936",
      x"aea26f0aa9c2d376ae6ed624a5858bf8f2d96f2b53e2e251fb835446d90dead1",
      x"37d05bf3d9a7993097721651b3e0d08839bce6cc30f4824a735d27bba75c2669",
      x"50ae726e5b09de810355aa29dccab19ea37778cc964919e232ae9d021ece95af",
      x"70fafca75d9155924c5ce61c6ab38c3eb0358efd45047d172dc1a8fa325595a0",
      x"e1cc9ff5ba7bcbe10fc7e3d8218f86ad164ebff5ae02a07faf0b7292f7844632",
      x"ce74affdb7aa93f6ceadab8ba35e1fc273d71e8cb2b7a6de0d6a25646455daec",
      x"4e16d49970b980d2cc60291b9ce01b4a47c401cb5230d22b3489d6fb43b3dec1",
      x"0c7a0a0604acc99cc24090c8ec54d7cb6dc0e6e4855e386d5e262f2f40412b15",
      x"7ee73a6e02ef382aff1d0275338d513b016b3492201c9b9923046503125f07d2",
      x"e2decc82ca4b299c978df9f0ba13d2980c977c806788ce3543f5cbef9126eb11",
      x"4d3247b7943e3052b5191b6a1744888f230665d774865112b290b4dd244eaac2",
      x"c6c40f7167737ffdafd051e76eb2fe37dc660553d4bb84c448f7f0b55064e5f6",
      x"8655be99217845d233e692c27b25d193cb28eb8a800784ba3b4c4b5e4dc764e0",
      x"26a5595bcca76800ab2dac45a00edb1c67963e4dab7048af3aee02cedea62d4a"
    ),
    (
      x"97d1e377936e28d1b91993da1f2cf97b63b334f86faca9973828f84279ddfb7e",
      x"cfd7d3c8527ddc6b124d47dfcb496f07806aa904bb068f79a29123cc97cdfd24",
      x"223dfa375074a886aa174866d3401a958264a09762b45fa76ea3403bf2556474",
      x"6fe41cff8aa3fd6ae8841a1c9f674cac0a46adc94ab3f4eb0b1416134ad43645",
      x"c2700e4b99d9489ad68c4ea6a4f6699a3a7c33e139827304f6010824719f8ca6",
      x"c96673face26a1eecdcae12081d07b710ca368e074236480be4dfae9e3303f81",
      x"0fe4d5263605147a80badb6b14f89d74ac2853b8a8b805fd095b4d88ca28eaa1",
      x"22dbc0be10f8c9195c862bf177c8fb0e89ff386c704d7bb72f242bd7121cf2ec",
      x"8d46a3c17b133c52ca52fec18eab8b29edc481faae50431165497b2f0b83ecbb",
      x"545e16649e92dc15885a099c5ef69ca7a717c0eed2d7dcc3a35647cf2e2403cc",
      x"50a5f3c49884fa95f904aaeba9e52144a2439abc7b7284b4a12d93095189b751",
      x"6b66f5b4e8b4f6f5d27027e605b3443bf55b3d89a8d884bbeee0e95557c456a3",
      x"82099103f4b60c0fc5daf618e0a9bd53a37c95945e6b3a49fb2e131462928bdc",
      x"743f2819951cd2bd420dc96602666ca692996d3ec249ddda36ff895ef17b53c9",
      x"e870fa3cc8e45536e2476295bc4309853574f09264d7876548d960701d6e9503",
      x"24e36c0c9090f98ccf65e96d6b596465682a0c09a4e11fe237795e1bf741b1bd",
      x"cd10ff3ca0cb1b21fbc6cb7fc47806b734961c975893431c47bd509a8ee79633",
      x"808e3086ccd2a482b91cce9089365fa60e7837a0a032b65d40525c5f5926801e",
      x"6fb105561a41d5f6557b425e6cc17c53c84ba0763ef226e65748fdf3712324c2",
      x"126c4ff0233b20081ca40f64c6c12d14e31197f7b3cd25664be063af73a56c94",
      x"bc56f26f5e91cdc51e0d39f40ecebcede48dc3f63e9d373f0ec0df298e0ff5df",
      x"abda03d8b9f08048696499ece95266163e32090befc6f772947e519f6ba8fd5a",
      x"a2b232d29c3d2c9fbc1c16588844a417f1cf91a07ab517e4052ef9a35e298311",
      x"bf70d3a8cdff42cd97a6570634cdb7c639d85dc3f10d047a99fd4940b9d915ee",
      x"700ec9d801566378c002844d7ea3b839ff215852c513c6c9e90e341359d70ec7",
      x"c1b64e12a9e0f0ba38f1ddc27ba9651db3ffaa62448780044d42cf9caed0324d",
      x"acc22c786e7b8db47f02c7d8f7026fba1f09d2c0c3da99ceac170c52be149144",
      x"2633b09c978f16223f0ddb2baf9baff0af89d4888379dcfe3756e0f2db4c9174",
      x"058626e3329608f51d0d645a35f122251b77e8eeb3325ad2efed2e6264e0d84d",
      x"04cab0c8392413e29b7009d8b4f3a5d51c46da451119da37d1c4a1f0755c7ec0",
      x"35dfc116266a9a07a02b99dc158df461c1ae5894c2dbc3bf6b34601b6ba0ce05",
      x"1a34e2b15d50dcada42e9d4f53a1db902a0382ba88aaf4031cbf80e0adf44e5d",
      x"2a59b7ac5f38d9b7b6b3fcc43de292dc38d6f4b25c09b3d0a129bfc0891b5ac1",
      x"113d3e4adc54f9a26501ef64b5bab13e26de0dcad06efcba40e4c8bc47463ffc",
      x"0ed695415c306d1ff8af346bd4d8d3e536828f298bdc85843e8c92cc601d92bd",
      x"132904315a03b6ee0fc629b35113fc1b9b2c9d939a103e82f29985da86eb4ac7",
      x"11d1dcb6331e7cb919830846bbade67d54a258f156d3eade703e2b001953cda7",
      x"df679d458600c815dbee39da08ca11311cd922bb6c326f01d7e498d6d67bdeeb",
      x"39b0b9c1b0bdff82b31a056b540f45ef34cc7f74b1cb2ac6c32be827d0475b9d",
      x"6a16881a2ffc0fe4855f454d7606b2c028ea29068a3896407010c8da1c0f6de9",
      x"6308469fe5498c1c109b9caff5c202f09933ad8bdcbc6266604292959402033d",
      x"a95df227569d9a825cb318e2d6adfd29d31850b97f308120aefd986a8e4a839b",
      x"1e54d8fcc51a101b52f10ac1a6443fc56293bac98d0f073109616b844c8a122d",
      x"b17df267c8a489c6bf5d1c2c71c1777503b728d078a600a4f6254b57fa63bf32",
      x"9452470be1325ce47f979b4186f0b4634d7acf14bf24ee213789c203e277afd5",
      x"3476e9f7a5a2ce55051db470b7e6d76318f4ccf03231f4e8d9a3f6c120b52b9f",
      x"97a9735f7190c06b7eb062ea4ac7cda6d00b67268eadcd67e3a07d7042846421",
      x"d347b7c13223075ea95759dfe99de29d391038d58971d3d34cd36a4196f6f1f5",
      x"f26a669bec9ac689309cac38a9c4ac23e5c453650ad872fe97b8416ccbf1a1b7",
      x"8ba00bd22a3f43bc2e0e0badbe9d2c079d6e9eb3c84c21fc4a43628f2a1fb9a1",
      x"e6de65fd6f4bf8dba3b970a15daf7830ac0708c5e0ca0a7f3a2b27f63a5568d1",
      x"ec418d7ea4622fb3009af58f039122898556705a8f04a0702c61f15669294b69",
      x"9c853b2dd6dd204c2b70b8b37674e0d356d9e49ea1c0ff87d2b1555b63c93928",
      x"67c0392ee58fdc2e23646745cf51f3502446119fbab5747de3d6ef81c537d3c3",
      x"87908da78d84408363e607fb219c959b07ff1de9ec4f039dd9cdbd90dae7437e",
      x"d77b2a3b5cda4f9ce767dd79bd8bdab6f0d4c687c9733f965b854248e2524ff3",
      x"512ed6a2100780a81635a3a383d102f691c035089484b7a556d67d3e9bd7dcac",
      x"bcc346e786d307e9398edc00daff7aded41374dc1d22cc284f2ccb5408cfb129",
      x"faaebb8c0956234e143719df89f0f7d4a04dd1aa2362c7807a7658c41cadcb9a",
      x"9418ed43f109f7de3d0558a2bc8fac86168b099f7e4258afd0725341fb20f461",
      x"f0f7e5a28071adf7083891e2c541c8e7bbb7459791342fbf2ebdde3da9e5cbcd",
      x"dce57ea7a6be5eb2df9bfa29c366830d075134df1ccd6337255f5f2a4109cbae",
      x"90a6801a63964e21e8da38b12363eaff49fd276b655dea25f196ab2825e3a2cf",
      x"389bd2f30f11f494d02ed888bacdce66f4c6bfb3fa431ff3086e2a813cb5a216",
      x"cd4d6fcd0938145a27a2d11bf55e0554902d2f09624731cc4bc3f84c2dce0d11",
      x"ace820c107a336891174d9967ce6a5cb3643785a496f147c4f61976277f9959b",
      x"bffbebe5295b469bdf6431ef3f9b9a8d909556a0bba6a6aeaf459b5c062cab66",
      x"7a23a680ee97e9e6a164c0742d221ec5d44f1799f491221f2831a82ada81eedd",
      x"31fce15464a85b738c7ec834eda69e183f1896feeb00e3fdcd3bd4d3af66c58c",
      x"1c7d68a9c6cd05dfe51805a87c4b45b7bc737616d8a241c1de8ba7c7ba07b66a",
      x"24e1034e2205096987cdb18c6d36a80c7130c801687fb469b364153b67da3d02",
      x"aaff8fcfd8e633150753b0388a140d5849d05a62e27d3167a05eee0063f9b3d6",
      x"ff1bd710ce506c9591c3e2706ba3c1c9a07a932128f1572ce16561677c860799",
      x"8b63df25bce11fe7de502acbafb412eb6b90f7980537e39cdcd890abac2d7a6d",
      x"c0e8070df4037e5e83dd4c7c905330fa46fb337ede04b8311d7de9c4cb9b383a",
      x"f96a0bd1db6ce05943ad4d3ef77b2f521cf18d1cfec9d9ac1fd0271769afbd91",
      x"28e201f2adf54111f741218adc102aacf407427a401d09749584dc43e96d8114",
      x"0518e3b4202eadc99942092a052b3037b0a5c4fc08f4ceb6f25a22171f1b98df",
      x"0af56575177ff3303ce35261d89648773262f9847825819db3d88ec40d8858a6",
      x"2e24c4fce33b2790fabf6b0d1166c501e4dc2b84cde59585344135345ecd9dc3",
      x"5a723834de16982155b116d49e90bde1ded6a744f383eda9d569b57c430290b3",
      x"10f9ca2d973bdb4e5408dbbc880a159cdf7bc33ba8fee04434c3e451cd270342",
      x"c3670f5ac2d1ffed61d2bb1e36bb2fbca81719fb9544ee342c6e9b07e931cfec",
      x"6b40f2b8bf75067af6bf0367601a354c1e9afa24a7008645cac0b6c01582b10f",
      x"b5a1c6a6653cd64742eb941b5c57495fd1180629aee66566462a60fbff4907aa",
      x"4279c5d9c2cbd30375eaf7670d14dced8a9057082bfb559c22a884a95b2cb771",
      x"ed66491f2dc3f8f7daed9b10e8cb560264d66ec67309fa8dd1f0724f9550067e",
      x"2720a7741e0bfc652e6a7149d1829b67672ab718629fdf9cde9a44ddc2b09d30",
      x"9a36239c4213e0f6129bdcebedf2dd58a119ed063e257f74af4d0929eafe0371",
      x"52ce919eb2d2947b93de288a7c526ad5c7100c49a4ec670a754e07088a99ffab",
      x"7eb0774f15519265ea9a448192bfa521d99e4046ae7a802e76f4a2ed37b66005",
      x"74edb0e5421baa3bd9a687a8937bb5ec229a2f77cb5d607fa10bfaa92ad92caa",
      x"848618b0f78fef30735d23c82bb7f3522972f2ae071aea7b7b70b9da05645bc4",
      x"51dc1cf1f3e8af8c2a01c9e4ba5e1a1f430099871f9d9b2ab809e49f77283a7f",
      x"ee6f4dc11a705b5e9d8e6959e321e4b0865753a45bc5c5a9849255561f412eac",
      x"076ef267d5a2ddf798a535e38f3cbdafe8d9cfb51cf01c48dfd158ab8269b4e7",
      x"c570c388d98c5ae9fa4773a6103cbc7546ebac985819c6740d5c622423903ee5",
      x"8e36fea17ed10074bb9c4f6c797c4d1d42987934cd0ca682f1814833705aed48",
      x"c30071883b3bba7cfe1d5018d1125775ecee6653fe0ad90ca5827cbca9e079db",
      x"91509e80f97d16f6e4d249857a4b9d76e90aa88019a30a067d4b2d5034cdcbd1",
      x"17b24e966c55b8f49d3b9196f62b9f65e6062213bc0a27af2ca3fd26f7e5c75b",
      x"e4032485ae1d9f7f060bb905c15d9b20ae0b077b034569f1fe73b21c4506dd3c",
      x"be9192fcd9f5ab8e8bd8de0d8f6135bc0f458e13d584c0da664cedde9cc1c0ee",
      x"eaed77b610bdadd38d1d5a687a64c1635866a7c5dc4aa7d1cc0bd7b09d96fec3",
      x"939d5837ff2db76eeb168f6e6b188f394a4c9c498f8f3ab89088f7fb54be541d",
      x"2f41f766252c3d5d1bbff92afaf8e2e7c6e8b4b8c2e6653455886bbceeacbd99",
      x"72f316faae6306c65af4c0a725148bb793c9708e8721b556a1b08f944a8d5652",
      x"427e8bcce9f8c543751e9c374c62636a48a3a00e1dfbaf99c03d5756842cc04e",
      x"8f9811258436555bcdfc7dae1cf7997e4040dab36723ca87b218a702f150a29f",
      x"95c940ccf8bfe0c270ab839725719db6d06013aaed3efe1cd48e0b2904a97421",
      x"d037147c0942fcfdf41126e2fbdcc582c44846cf0c6a43bbfae350b1c3d17f2b",
      x"1f5088050ecb57a85851125679f2dbbb00b2f857ce18a21cd53506f186d0a8ad",
      x"06f434dead048b1326bc7cb179d3238db62005ecce0aa696b479d7fac17c9f71",
      x"8a5aa6db4ab2e7d0aefee81002bddcad4a25d95003e1f30606b6f5bb7cd1a48d",
      x"e3fa392bfe93bc5d56027dccf2f3a9e4ae1e765875739f40900821c8f15e4f7b",
      x"eda1eafd54e9f6a007578957e638a58cfb62be251c8a3d91aa1bd0e38a417693",
      x"91e5ca30500b35463d22576b02b9f9e00c32fe2be551800962f87b817299c105",
      x"f7347ec3597c416406a668c0a85eafb54dc24fd4b9b25ef67e63d1ea31e466f8",
      x"d614c55cca700ea847f1b64046a56cddb16f658b21dec31af689de10c86902ff",
      x"cbdd15e2713b4ed32a1f42beef415b5b4ea6187ec79f24f67517e7c4aa71beec",
      x"2aa7a8f7021c4be3fa330349871a7fc6f58dd99ace29c960da577c1a1eee286c",
      x"5241ccf144e3f01547c934927b54e90a4030f080cdffe5ea4a5082060c2579e3",
      x"6894e418f43d675b80d97997c320e3c914872cadc8b55e4eba53fd6730ea3c8c",
      x"3be525c20193716d04a93d5b9dbf73924f7fc24ee8baa5b69cd04cc5d9249dd2",
      x"1c26151c83a917c880f1b9e1cf3023deb9a830020d22803d33f4675f20411ed7",
      x"6544c1346c072b4ed1bc206d8f3575f4f76354dd5894e5c7a27807b4433309bd",
      x"2f694242209a1ea09176918af7aeeca38d8d28cc282e83ffe28d8c30000b40bc",
      x"ae073920ca8d657810f20c448b8f235767d1e9abe5531cf3ff36b3875fbefa2f",
      x"c0fece39293cbed649e27a264ea82f5fbe0954516c98c4d419a1f522ce310852",
      x"f551583727556f627e5060f39ce93c3765b78a3b15a6863afd9e3b4f5a4e63bf",
      x"d9f44a7e794feeeb864027529813305994087d0f2a909de5efde6acac83aaf3b",
      x"c07dea3d7e90e2b8c984515c43ccb2a98770c920cf0ec122cacdb7688ae8a7d6",
      x"520c61b3dbd8e9b35f9b1fc2d9b7051d8eb28cef8ef5c2b458ff46149538817b",
      x"516933f31223c25cf86b0288d75c18358b1c70f048310fe1dfbda917793b6ea5",
      x"965ce5ce5ee340e6b7b1d1f513817433dc3fcf0c2ab414c3edbbc1812c3580dc",
      x"e215eb11da0c940db023b718f208958b46cd1711fb8b53b48373171249c195c1",
      x"5dd6180fbe1fc04f260a2edad42a98c1f41a2a3694e8c6722a9c8fc252e6b92e",
      x"6767c9352b6549e0b6ae03b98895a6fba5d0d4d2397156d864d39491aedcbd64",
      x"e9708da98daa85c5cf91226178cbf1a4653c6543c6906209032c423db662266d",
      x"10a1570169119d611ce1d0dc69ee0ce4af8352f27e6bb9535b7dcc59aca0462d",
      x"e10cb21994b177dc587833cf8180bdcb33f0aa9b33b8aaef65a9eee61a7a911c",
      x"2d2392303028290b04fa21467a83581baea71a742934758123e390dafab2add0",
      x"628f118e097104e5ca9701b62c2f2c224e6b6a103c2d11d4f0e51525aad07e54",
      x"35f360f541cd2d442d2c2695b98505b5c995fb212b6828fa83165b386835218e",
      x"46549b97d2c7bf5df43da07b578248159037d6f68b701ca09a5fdb1c5aa0d1ae",
      x"bcba1facbc009786aaee1dcf932fde749a35772a1a4207d1abd37dc57add159a",
      x"66013891c17393557b058693201d6f4c5a3cdaf61c28c0b78053a7cbc56a1cec",
      x"60734870c03a84557503e72caa9c5b833125c04d67f2f6ef23446d8d5f1c8e71",
      x"ffa3824b44ce8788d77e0a09067b59bfc3fe8aedab1853c9b063a19ace4b839f",
      x"218c831d5189fdcb6c25c6417a1ceb65bf59f5ad340cb9ec1cd69d4a5df32dc5",
      x"3c118aed3447552552eb91479581e718c53f2c8a7d1d99b15a99dfc961532d97",
      x"2a43ec8b3f5ccbbae2d287b5014218ae7a65f65e71cff78c4a1a6ad283c47d77",
      x"789a506faf7f0e8e6d9af72e5209f490bafa8918a86590a6e5c809065019ae45",
      x"ce877a5ab4c278f20f660f080db3e4084210415ee0a1e99c3664c9209887eeef",
      x"91730bab94463ed3a288506079a0b59e32dd6858d2ac53e3e10917d78432b1eb",
      x"cdf98ddc2c5483182cf68a3eb25bc98561c24f0e8425e263d9dc2ebd8911bd3b",
      x"95380633b5ca544d61a9c9deb34a58121fd0fe32c29b3cd95905708b5ef551f5",
      x"346d1d5467c5e23f543c3e7a73f833c9caadcb5c440618b671d9a2dc5a000ced",
      x"c7f40d2307c34043f5cf2fccc0c9c46184259c9c4003a7885d7e68ade17edbf6",
      x"e8369e2f5ca2fd6f1bf085723859e1da299d3c9f9fa0e5d078d64904b1a8009a",
      x"c3804db966e6f0ba4c033df975b9c73ebd7ff1f288fa0ca7f844c66b957359d0",
      x"60cb7ef2561192540b586bc914a8e073047b1dceef0748392ebe2375091e6e92",
      x"2dad2d063d8107f8c46d80c92e56c0edd6fcdba4f7daf56920b20eee48b69833",
      x"e4b1f0a8585af2383f2f25d8558fe10cd7eb294e37c5ae96c1c8f4d8c8cdce48",
      x"1ba62479e17122994d43810f9e3335c85ae8046ae1d02662756c2bb5344674ba",
      x"80e94a4959c11baee63a535cd2cc6107b9e658025ab4a148f8f738a368f4a436",
      x"e55102a5d80add4ddcbac3b333f8a698b4c31a31d8acbb5d02c673d425192c66",
      x"13b5b683b13c863e8b1a44d273ffb4b5265b76368b89d757a10d53210a87fbc8",
      x"d7729fb9e2a16d0e72b2ef00abeacd796c2e4cd48dc13903f0a2a7dde37c86c7",
      x"f562384dbd35ae15b8f325d8b36516737cd5668c90cf5756c1a2b236fb87ee93",
      x"cd8bf2d34410a2ceebacba16cb080e8ffcaead7108d4403cf15cd1671d3c840f",
      x"936f8bca022cf118cf0f15a99ef8542437ef4f9ea1f7092247ba055579e1a941",
      x"80a20ec5e1ed72406f0fc905aa31f81f4f50f363872d0f3e607e2670825a6daa",
      x"84e01d296fe51fdd44051b03cf03f9412e24780ad271855cf0cd5440d99bf8f2",
      x"2c744389dfbfdda9fbe6645dfef29c339dd4733835c1501d523d46a79e620ed6",
      x"6f53ba59a363b0e0c1529424a61dfd59c4b019796a28e6f24dc5fbe92336cc96",
      x"d82b65ec1dfc42001a571abfc76f65232ace3b859e7be63cf1aab6d2ca1324be",
      x"8fe166a1509234f0d9bd3ecf51b454898e339dbd9704dcf9d430b5657def3659",
      x"0398dc52e46538429371fc6f3305cc34f39d3b29034e2604bb5624c48134607a",
      x"a762c4dad6bcd586600966f4c83243113419b63b9c133149731a816a5928722f",
      x"bab7076237c11a98e3ae23a9e4c283ce11e6793234a3f2e7bded56f153d25c33",
      x"cad9e2eaf823c5d5009966d622c1ff6ef72ec936be8ad90234034c4dddacf4c9",
      x"1c9fa3e2e1ef75fcd405138b65c24a8acdf6bf37ae8e3ffa2185de20e43e3aaf",
      x"87d18e33036cb80c3087c7a45e594f56f8cdda339d619f3491077a95ea82b646",
      x"cd3db6ab1d88e7e3b0d8a9a2f5dd8661312bb9e4b6efea0bda911ba4183527b3",
      x"4f182adc5b21321fae69a113b35ce511c4ac37e782aa3bc5b0a11c8d7138f709",
      x"1d9e789fb133daee92dbc57c9963dae4d1ab2c3c52b1007b13f4094b90840b81",
      x"01525b6fb6d36ee251c49bca644a6bd7e5c2f14c1f84b7a6262423c170cd5420",
      x"cb1d39d39bb675933d6d806534335bd035230b47e61412264694fc1e833dbeb3",
      x"2b3e1664076105e537ef0421357dfb506e6831476e58248d37e4c74321e9b095",
      x"ca1a833b82f281bce147d14475ea21ab7699abb08864f3ef435030b2bcece651",
      x"2b798055f7330afe6599e3adc34e32cae94cda796dd7bd30ef8274fe969a2fc9",
      x"0812920da569ad3f9aa60c9eef9f3c4cf26746424923ff99ac869123cd2b0af9",
      x"4a924cc222f05f83f32f32b6b3f763f9ef9be580b5120a149a4a7c366fb6b235",
      x"5b64b57baae28ad6ae9164191bc08a0e8dbd9617553b9e2742a2db66c322d75b",
      x"ded34903f72d5cf5e9773333d4176466b30dd48b16ffcdf8066782b7c84b26e1",
      x"13d944a3dbc1e10747e4bf596093e92d07431483fd1bfbba11e400aea1e188d4",
      x"6b528d31c11385e05a6b0003739c6be2bd7fd8133a688624dbb63780141e7546",
      x"380a0238d571c82904789280806ef92403de4a43df4fed6b8945f6262bf93743",
      x"4b4689aa9a23ceeb272e90b2bc7c664a8dd22a1da09cc524dc86d7eb08211d44",
      x"23a787b5c94becc5d205d8677ca14d3f3f0b9a882e3729d4d2b7f7a2f9a2d568",
      x"3fe01d83cded24475be7fe6adb5d58989415a3c3bf28861466db732ed8cec554",
      x"a19942f17b53f8d0453ef56d0f6c83d095c3e75d0fe23de80d042181013053d0",
      x"122b7ca8ffed2e2a916f0ae7d3c36315e92fa84187bd4f6b940c8f5a3ba88cc1",
      x"de920b221019d5445ee6aeeb877dbb26a11da6a4d060392c424ff3e1013892f6",
      x"ee17b1c74e299b23392107eb677a4dcc2c68ef63b8b846cd4f5dbdeb1fa8b41c",
      x"cfef823e53acfe42c6319cdbecf4c68d5d7cdfe659589501d4df51d7bfd549a5",
      x"0b5ec199fde32bc2df8f1d115e729bb172938aaca73328ab8012ab16186b481f",
      x"472cb293c9476c267d5b252cf097726080cecc701d9f9e294e7ba49753fa5ff3",
      x"8476b6646105f1b49f9b68d3bcba97e5826f8f100071e3e2b6c7b826d6fa9a15",
      x"84818187d151500e93656fd5d41554705e6169f0ba97f1c7b2d168eab5d4ab81",
      x"2fe617d6bf423e79c7bb334fb98a4b2f26ae7ba79971212cd5a9d1739d74adcd",
      x"482eaed0a481f99c6bef418ac52b96798440d7e070df4ada4d623792bc01426c",
      x"402a71244932b3d48547638babad2526399adbd41015cd72d15688580b270edf",
      x"1e8cd1c630e29bd7de7d170823186cf5bd390f5a968b3369bbc89f162fa92cc4",
      x"5318c820826bc259518b54aae48c22083891f1077a886be2c8784c509b831082",
      x"b32e7a44493bfa3c9e3f66cf510c6ca54acbffed0f80e22e57a5fae78b79f2e9",
      x"63c8b547ececa8bf37896dd2a5c719c69f73954bca0f720c47a79042bf53a7f6",
      x"e47fd6468d5213bf30ce3fc1071fd9d559942819852cd627dd892ce5af887f4d",
      x"481382bca310acf8cb15aee88d0732bf5447fc65d862db085ca1addd0e305d89",
      x"dbc54e1d6e4d1976b1c93ac389df816e033e26290b9cf12bcb9418134d88e033",
      x"0a1a606e26300545a57da75b76439386c4239869c42490ce73d1dd5d827e0f95",
      x"81114e9fc5494f470d4d98943ea49ac2c41ec502af0c7fbe04f183360c0b9ed8",
      x"0048c93002e9e22576af74e6ed5480d69558d019f4d013b5bdc6158ecaddb5a4",
      x"a67019c59e5853cd07fe55de028e686f24ff6d13f45ea94225892cb3b5af24b5",
      x"842b6770a0cd8d004878f177d0b0c83a5ce26d2625eb33160772436de0654e80",
      x"3aea1ce30c4af649bd47131439314ceb5f525253b6b18c5d17e5c8485715a347",
      x"e6d108323726b3ae58ee1ceba6a9816ca2f7609cb27e3c0bf4a4e13d9df52b23",
      x"672cee35b7a34705f53436a7df1169b151cbfe552c46d3cf77119d7766c3315d",
      x"3cc72fab4222144230bd1c1072ca02a222406e588a0bb62c16d325d98e42e577",
      x"47d959cdbd376f7c5d77c5065ccf6322ae72a2fcc5074b7ddf212d97c8a3fadf",
      x"cf868e34b9de76a68743cab90de9d7e8cc90faf4238c37dd67c5fbb2fbb0895a",
      x"c6a1f5be45c0f48d8f112476125ba5ec2f30e6a768c89a9b1c487734d5d4f10f",
      x"242a146719a7f97fdec9e6ac441e13b243bb0bf00f478c0027db8b15e0c6ddee",
      x"3af1c6f754285e15076e293f42babee8e4518639b4d7490531749248ba040f5a",
      x"c6c18b7dc5749a16837c090389aaf56d3beada1b31d74ee748bbaf034c90cd8f",
      x"d8c4cd7eb286928691f64fdd7a0cfb958160d99f8220ad68db845353506f06e4",
      x"153c90b51c3a766621387e2f81da67ea6c77988af9c78c1cc4ed465170841b07",
      x"d72a260c35d872ce8e47f3e4d506cd1bf85c3f34385a1693b2ecc8ad3a36f699",
      x"fefc76e987ca41e925996b19c407b31699c021c71aa3e297658dd8ee03912176",
      x"77327ca80026bc5fbac9330ed1e24212569d40ee2cf917eb40589f161313d23c",
      x"6611b13d38dfdb4f4133424e98f5334c4a4663656c82f7aba023fdf72442a372",
      x"986c879834962b020a7c0125e165a3f79c0b230efd4f1e7a88c878d7b1c6da6c",
      x"533b75c56e0f5ff66704f9cd5a1271c5a1bec5c82492747bec54cb9d948a3fd3",
      x"0086c56dffba5b8c6872dceba8cc948fba687854a590567708b3a992433a7088",
      x"f19ea699503aab35921ffc5f831cc4649b16151cfe9091050c5ecac355e6e5d8",
      x"38a9d396947403d4d5fab6b1c4f2f16930f76774d7b476ca48dbf378e59000f9",
      x"8a484decad4db0972dac7a864af5f96049fa64316dc57a9f89d74334e9a3b35f",
      x"2edf055b72f054504f55f07b3dc3ac2938187208514d4800a63815cd087ab38f",
      x"d2c5137ae7a671373bb8ffcd3f6174be8bf748266cd104f3b34b922a97494aff",
      x"4b22f272343352895c32db68425aafa24224090766a7fa0ae4d9d428ea6117f1",
      x"2635302473b08495746456c252588e838e68af64c03d50bb663e7331006c299a",
      x"dd527182651083a9a791caf811bff43ecb864d04cbfff610f3e7d5e1e4746ca9",
      x"01b546b356de31f481c5294d7d0d01eef7037a289f517a334c269775901c157f",
      x"331a3b74141c1bfa12974cbe8968389e330d4ffae61a6c6eff4d3eac38d65aec",
      x"c52de8a0eabbb8ab84493cc11c2c04b1d1a3a4ba318d113a1bb601fdcc392361"
    ),
    (
      x"8841c11b27dd02512ec65d4d86487dad56997280f061a083f0e1163f93c4efc9",
      x"c7110359ad2d256e2c757ddc366d9acce1c37f3fe81c131b6c442db4839c8655",
      x"f746d5ec6e03627052a207881feba0f992f07f3bd1cb895484eefb7d2df0c203",
      x"115c2a162f2b655f7a309c35116f97a2eac7130b3c4355a3a248f1b2c3723451",
      x"f4be2e41db107919934abb12af37cb2ecb508172a1fad437782d0cfa508000bf",
      x"74c624792613af4a31f658c7785163d3b6949e15f2b28cff34e96334c6d4a72a",
      x"0b2c622c36a3a5cfde9d9818ddea8b93bee2a86635778bd58232e531bc5db601",
      x"3f67f2d9b083176e1b388f477335a32e17c47423a873bd7f6085ce865d4e329c",
      x"d1e870867fc451f3286cbc2a61ac40945d938c02dc040758a2073eb6cc877692",
      x"ff35458d01d970b0c64803b1f2a0764db3d94c21eb4ce59de143748abb600396",
      x"67bedf3dc90c7a12a4ccda43caea20367b19707f3ac72c89777dca2c66c6f051",
      x"7938a87594c4732ebebfd1540d819eac47da98704a8534f36d8d03a7584f763c",
      x"5837ebb33048dbded1b98234fdd797f39a8394cc94128ac1f763682d6e31eccc",
      x"6c7211abd8d5c9aacaf2a90824977860a66bc1b615fd7e32692f21f5920d5860",
      x"f43add76707947c36592f61abba0be66fb5d3b005e73d3d69af607a13d5eba9f",
      x"aeadb36be96647850ee65fe1eeed84b92998d638592a84f23bcdf24a300b9250",
      x"e91364fe93369c7112d65f27c3cc78ac75feccbd6ade4724761c692d8fa33cdf",
      x"a686ad66801a6d6d3e396726bb8ad4b4308b7526c31520e3efd6872fbce156c7",
      x"df282df165a6cd2b2a250f04e47e13f44bd313c4b5ac0a6aebf99b2a37814fe3",
      x"b1f92e90f83e779266c578d53e08137bf736315d588ad9a0fceea3d78a9ea39a",
      x"03370d2be65e866833ddf5952e3ace7764c3aa14ac436daee776c57d80755808",
      x"16261069da5f8ccafd896a5b02130f7c33ea9f66bcb28e9d23d10aa14e6deb01",
      x"4622fb36e82540e354952f6679aa8283bfb0f66ac91e34824d0d3ef045f66f6c",
      x"641f1344452607fc2b223a180cc1277a935b427e1c24e44f213aebc0e7176c92",
      x"f6d20b1b55aee10a63bc3ee8e02873346ebff51545b6d34b641f948c5cd52c45",
      x"d9ded183428b7fedad9a45a1591d19cbb6c3d08e16efa90b8144260584bee286",
      x"576c7f7d2d1b74f5bf9c508ded58142553b2a850500728eedec16b38630e8cca",
      x"d40faf4360001149d9aeeedbdf4c65e1a9654a74149af805fa6f888d12d78494",
      x"30fa636b40cca76b927a7df724b019dfb1de8d859450ebb30c5d6560143c38db",
      x"6299d29b183c37d42a88f51bdb02022a9a7719828569f6450c73d2a2f817a533",
      x"b103d3ad9a6c30eee97fb2961bbd50fbf7db28d6eb4e6b1f19d3e9c45b2e12d9",
      x"92e5cc4799b83fb6cfb9edceb1442c6b3f117e66608722c26d756ac50df8f35a",
      x"8b0ad2c7d28571da3997c6ab883185f91c6b68e3521652bf7640758d10d4d57c",
      x"e730bb41b29abd1c5a902b7f5e9389bec6be41e83f0f0bcdf5f34e80084ddb41",
      x"94eef35bb0b0275a8c16c557258dc8cdfd27d041fbe6658bf4c41a989b81f97f",
      x"f9d52e772af00b486160940278c657e7305aa1bcd220610f1c8580be211b9caf",
      x"6cd22f45a537c45f3c9c9c37931ed6e9e51a4750cd35e57f39127d8549ac07d8",
      x"0fa13ae437cd924de6880814fad0c1e04c99bc19ad85e5d8850f6cd321f74eb1",
      x"5e4ba5163e50790f383fd1686d79bc150020b64c51191dfed24994cc75686890",
      x"d04ae00d61fa803ae08086f3fb126db0103259c16d1def74c7bce31978b9816a",
      x"a4592a63cf860daf9e4ae9eec8a09e197e4f8333ed166c747a5df21d01f5d9e5",
      x"ea5e26bb2af3c56382c3beebdf93cb0cbef9b257a07c8ea61130b960af63e24d",
      x"5eb83a49dd6580269be2bb04cadd795f8d2ecdfa629e6d38cd1d4dfc87655007",
      x"3ea9148ef00f7e81b041b77f6f78191bc616b017348f5c7314faf243e2265959",
      x"919c13f2964f7fbbd35aec4af9d6cb8e7da108dba797c3229f38fab9e65f8f82",
      x"37f9afbcd36fadeaa43f4541bf9cd7f20d41d0bfc3d05ae33b8eb43e3579f7bf",
      x"086d8aefb08e547f1d1fc06a6968f2ba5d21487bc7293b0cba4e41faa35e44af",
      x"fd0ce0f38a7b8c780361aafd25c25595bd4416bbace5926f944d0a1aa70cbefc",
      x"ccb2b3865317acf5d0dc4c2c52db8ffb75e4e645b233b6654fca559cecc6a999",
      x"06d9618fe12f6216ef94a094fa40ff793283d228bac2b25fddd29bbefc2c446a",
      x"dca61d44763a9c142f3bcfa7b4f7806b52d5361ad16a2fe8fc33533fe0b4c63f",
      x"9350e7f5bc9409727dfd09db3e315ed226e1544c8422e2183c2ea4551db61f3d",
      x"8495673d0cc8afa6f91358e96d4055c9dbbd6e1e2adcf275fb38e4a389d4ecc1",
      x"e64cca19019fbc4835761a8bbf00a405326a2153ddfbb0b898d9b4b45d971e56",
      x"fa4abba5dbdbe9cfda8af09afd7e89c6eef715ce80f459e5d60d772ef5b27789",
      x"bc5d070a13716a1259306a6f65b3f9e19f4cdea7d69b2d5d47608e9b8f085768",
      x"d90a65cdb3a80f71d62681c12f3413dd2fe8224c2a2feabbebf54ee9230311e1",
      x"c03d64727dedde09375066ebcf0700200fa201a4a7b37cd5249e8be8fb535f45",
      x"5ccccd56ccf6449df53a78528156ba56a52306354fc5c2b39b62c3c60a200846",
      x"8bddc901e027287791d0c8618270390798ecf9b682b8bc48cae9276c20e29f66",
      x"ed6ebb33d82dbdd633dbb800543d471c6eec2dd82c8cfc99f416bb89a4b57ec1",
      x"ae3cb515c259fcb2f0f4194b24dd55397858562f627a15ea4e249674d86f4df1",
      x"744de72f03a2f79f846671fa8fe4d2a7dbf2595db4100adad5bf20ff44eeaf89",
      x"e713245726e8d5923bad3390ad65760512c70e079c561fe6870aa957407044ee",
      x"7489667b22bd3ce3becc2c7d024c1cd871af8ded6cdd01a73255bd0b20688b9e",
      x"7291190b127e087dee4adcf23e10496d1e00e617ee9b73f685abc749321e8a04",
      x"e909622e6405ba5c6ce1ba4232a888511784c3e6df93da92914fffcee2e93ba2",
      x"41bfb9a0ce812565de6a115b21e53a2fbc689be70a1853c0f106ba9f1de7d9a8",
      x"9858839ad4ec0b8b5f41965958c2eb55ebb5b0ba1c0acc492421fb4ddd38b3f1",
      x"d15b89c01e3e6939adf01f4dde3ff082dd8d48bc1466a750123eaf0fbd416ca8",
      x"606048d8b971dc645de46999c4c03dfea41788ec83d2c96946fb23bc656cebab",
      x"8121e94543bac48e7b5bf6eb97be18da1088d81dbe45178b775af2b959ce5f32",
      x"fd9e7c9fe26da5ccda65c179ea1e105aac48f2b6e2895a3a546edf77f74ef7ac",
      x"25b67e4ca96422575a0729593d2652934cfdb2f036ae294e2d118206840b0c14",
      x"9de88a094656e8cdb2461ad00806a944e6ba255a38d27fd02c4681322a4a2847",
      x"a0391afa9b103de2f9ed2d7a88a872c38be507645743bcd70a1a87b869fdb836",
      x"4ce2e19f203dae7f17cee3e503485f7e42e267cb761cbc36950002625afe87dc",
      x"e7e80459d9b3cd4a4d58fe37fe59278b3f8854635803794249681d39a4e391c6",
      x"02c2aa480e04c76ff7ae5c258b8e52884d8512852468cfc9769c75eb1a83451a",
      x"d0588afc03982148583f372c993cc0e5df922f6f1a403a5211a52a1abb5f44ca",
      x"c9a75c7ff6dc209ccbf7b3556f5506709e737078c1738bc0bb71d4ef1ec89464",
      x"d53ce87bd3bea85f5e662d1c6e4abf56f0ab0b66289c573c2ed45dc6e53f4352",
      x"cd7eb40b07341d6cd40584be18f26099a4ab45de97dd77455e3a1b3f1dcfdbfb",
      x"3411930abd456c60f04c5b90082ccc6aea51d6870685c7e20acbc61fd30ae8ee",
      x"31002ea4fa076f70f1f0e49638af949f30c5e30b21cd73afa3968724e0fb786d",
      x"d5a33b74425cd7d7eb0b7d90831f4e2b0537fcea0b1a1f3d9c96c918734f6503",
      x"71fa5eecba310233de29bf1b5f9db3031bcb2b372d7f8298a63770b4ee459aa4",
      x"8c5984b1352cb270f5979caea847eae69e2753d3725ac129436d690ef9a070c6",
      x"23818e20721d0fcf4988e0ef5e1fcb71fd09c07f6d2fd749e041ae00a780adb6",
      x"2ff0f08b1551e4dd9b0330966a99f18a87ef5cedf47a9175150d886a9c1711c0",
      x"bb1b7db0700adadb68e9cdb290391292da0e5310551fecc7fc42bd4e96902b70",
      x"2be9deb918e64c6dcd7270d32ce7850e4e3a159cfd89787452c14a9441cb003d",
      x"38f87bc8f3116a0e5e3df54c4eef79c599654a6b38f7124c2695af485fdc255b",
      x"7259b2ae772c0c73e0343eca1c9e8f47105350bfc45e8aa687e2f731a8735c49",
      x"1f6b1da907a613e96eb0fed639a964493b6b5720a65e0b7daa6d64eed0f7b115",
      x"5996d0f4271c072ce425d034e108f9d18fbc3460236d369beddc2dc9b4ad60e5",
      x"96e4a0fbe3bf3edd8c1d99ed73a0eda1dd55fc5dabfe1e8727d1df02c876ea19",
      x"1ffb8c2371f93f44ef505d7128088d5493bb616b33ccfecf4f34a7716abce1f5",
      x"a49901f53d68194908c6b1b59aa43b22c6814e058bf72320a3217b3fbe55d32c",
      x"0ee4b4e2f43b0cb42cb75561f01c0debd073edc70d76d86cebf5aa5a625028c7",
      x"7f15ec705b9c02ad43d8665491276a28d7e81ddf5a5b79e2abe56a1ce89d7083",
      x"0a2317d2cb04d4befb78573ef3b130108aedf7a375c0583a613632ea39b99f12",
      x"7417a4b94d29165c590ca9a6b8d720c764ee4abdca1c48ef76062322f772241c",
      x"9a07e00fbcdb2150fcb06f69022313c1b61266440a30fbd62f12079115fc3e83",
      x"2f7c614297734879339b708dfcdd654837fe38e227e168d934fa31ba9e2c8ac4",
      x"d253fed546ab1b2eb51af87f1ce16724615ab3a821fd0812cb5d0fbe848df1dd",
      x"9ddecb2810e9c6ef6d40937fc2faef1f24227292a7608a3daebcff921d52b0c1",
      x"f1e641ba5674f7694f5598e07b268081f743958bbcd0c8f554988bc0dc2c993e",
      x"ff04fc67f7429a41eb6eebe2e6f1987a09d728b9b6294e42769ab6b3a61c6040",
      x"d944bb76645daf236f89acd954122e3258832401c121f7f5bfa29d6434e474e5",
      x"cc4dc760f53ba52737d3782bc9e9f8bf52245d0ba4006ebe12fb247661ed0954",
      x"7ee944f62b4d6518f2c1d38b45b0e495ec2418d4c21294b2d0c32319b9b095af",
      x"70307dc9f755de4b7adcf2bea9b541b21b7509b485b8a1ef98f8287478e6f129",
      x"599986202fa57baab612a8c9434717be4f3d3a7df1c3559f4e87c70cea15724e",
      x"a8277a215631d5d8da2582c984979cfb6b387f20199ac78f544c217fb3819bf0",
      x"323d196541708abee99f4575941cd100700a564ade323e29f1031f1c4443e384",
      x"19d527eef1d9e6593d6176ef2105c031f5533a89826de619326c4cd53d91b45e",
      x"38610f1fd8a7a992207e447b60d13672493255fa1bcae5131ca03e4ea9adc8f1",
      x"2e164a07145726998eae1c5fc83ad3e424241d53b9e806a400b317beba14e9b2",
      x"fe1d6f3f743c3be73e9f1fd2684e530b63c40a165d4c4d5415953e713797ff9a",
      x"f1c932011e1a10d548afb48a64a7c2dd9ea709dedce8473239415f7f02ab20cc",
      x"ea9d74e26c37e9511265491d1be47e92109cebea038fcefd700f1cf538092d9c",
      x"09adc01d6ae95bb5b9adc873bd2b60b34a8c1f2515742a384af0f54abd3d9ca7",
      x"31f239082dd27ef51a70d625916f3f12f0174f246a21b6fff52697895147c87b",
      x"1bf9e4d8319092c7012541081101a523492506ac9249f4c019ee00f61c109676",
      x"aea6cd37cc84111dfb73006ad98803abfe4ddf85654d388589b49df69f841542",
      x"835e7abdc3c502001f9bdd6fe82d9073ab59ca0839c861da56101cbb519de7f2",
      x"18b4b15ae85f9ae42abddb45f233a2e86c1f0c8d85aba3821f9b2edbce776742",
      x"45c6ee234b899eb3b0f389d653c4f531f4ff83978dc1a011616691f131a0dcac",
      x"d6a8ca31b92a27159c139e0e39e0cb47964c0e27a6685c7cfc13b2221935288f",
      x"9dfb3b36a5694128b81c7be97a60c50a3219a6b7c2f12230ef417e08a19e0f90",
      x"afc80e0f44dcce79b8126d6793dbc4f8e0de221eb532af415a70c48318e94e96",
      x"754291b7fddc544c02658a319e07a9700c9fe604f3decf799da92c8ddfdcbf45",
      x"6fbe6e383c58c9d376282615fa42c726d587431fe226de074a1a26bd33f28544",
      x"e487805e821bc27497a491bef0baea8c986bfad87f77073bff6cbc11b76bca54",
      x"78126a074cc4bcec4ad9a7b49dc0aaa78db3f2e692d0c830fce75790b6009f05",
      x"f232853ddce65ce04205c86ff2698be422d09caa349e46a435a82c8609627e85",
      x"d188472aee0c5bccfc712e6b979209d151feb62e4ca21a8329beb0ea8a64c600",
      x"44dcf58c02da0bf81efa16cfac0edc3182054cc7f11d35b56f8da71449d4c436",
      x"3041bad7fec27c673d50b6f369879b8983fb580f1434ba118e8eb4451e692f3c",
      x"d966d7887ea38c1df665654411678b3b714eac6917dbcbc68eb3310134f43adc",
      x"4de59dee1734f2954418d45030a9d641c0623a3225ca7c40fdf7838c91d19744",
      x"bfb92cce1977d8bad14b5ef1df0e6b89732e35989681269865c58010959b1c8d",
      x"11a60b967197f25b62e1fdfc85cb0b96daefe39e7ae3183116622b9a6c078ecc",
      x"e71c3083629ec8a7fe283f02fb259ac40119ff5ca18c4ab0ae568c8959d7b49c",
      x"5940b9aeb20f89daebc384f20c6b9ded5e3bf2d47eafae8276e06c289e1dfa91",
      x"6095c50e7b8a1cdc91cbac497b1bd3de2d448a1f20d554ea4916e7d98f615fe1",
      x"a62a292cbb275e5ce871b359d56fed34720e943a1836c7bfa5149918791d575d",
      x"eade691c1851adfa75a3df639c433f96922b050d680744d0442061d178a9cc6b",
      x"bb5d820e9dd9f494bf53ef0d83e7cff19746bbffaabbf25072c6980f8dbbc287",
      x"7cf0b360afded5209ab82a33ae90c1cbdb0d359241f1245271146fef0fa79e70",
      x"f2d8ff363f28ef704d2b595033fa9f93e81c7cd048411786c36dca25c7619fc9",
      x"7f6bdb404defc10d6bd24e6be4a3b4a16da4301c67173f88f9b49bee84321a07",
      x"5a2ee0039bb243dca33eafff37f7f1b46f59a7514908d1c61a835bc104bc7f34",
      x"3b723bd857128f25c369aa810e13a509beb01d85aeeb0510a5b1ec70e83416d4",
      x"67454a4073acc1f59e28b3581b5db2c08a4f0d4a5a7c6d886c57b3f418fb73ff",
      x"904b0336cb4702ac0dcee4cdc47947e610b538aa0b830e98f1aef2d480f3d22b",
      x"bbc7e9f6b087fbe341372abed9270ed3c5bf3b74b2ef162d285e43811e815298",
      x"591457f05d10725e2b5e55f840e5fb5fe5ce2a5bc49ecfb506905ad325d7e456",
      x"fb6d40537057766a7288105fa08ebcec5e16d3c36d2d19afb1e66fae9351cfa0",
      x"3bcbbe4fa26075687a608692df58156900b6c7bbf0048b0af499aef632b5d35d",
      x"d321361b16a88c395af1ce55646ba4f694a4845862f9b5ec4f01ee8596bf70ec",
      x"a2eacc27b96069cbc95a3bb6f7db2b44627e1694bff574501b828d21a03a61ed",
      x"569ae8af6294877be4371f28ab5af3424681236c97bc8515163e7ffffcdfcf26",
      x"8c503220ce984fc1dcb648d2faec525a39c1b44d3ae27b5964e59574a62f2944",
      x"da8a263e4911b12b14c06c259c1579d6775f8aaac13986dd4fbf4954eb278995",
      x"1f8cbc3224ce94ecb7b892651dde586ce2fe4afb3d60cb4a1257ea589c5fb9da",
      x"244556de9f43f355f8ba92df2fbd71451a24dd38597280e3cdda83adc8b76a31",
      x"229582abff88f5ee0da9cef3fbc866752b505a4ebc4f74cf235ff457c45f0e52",
      x"955bce4dd44c1acbe25370fe18b37f39a773948684e6744b527182646a6bb39d",
      x"009878923ba2b962f7733379a711833bc62f37439224d30e786b00afc8edc55e",
      x"fd3b0519ce6c6f8f9f75708e12570e35a80ae98474076941c6398a355c798363",
      x"aa7bf4add8e74abad89c8f5d750235c438c2510784d64e85ba7ab614058a2506",
      x"8c5b54a9a2a0f3683c7d3f694287db0ec22b0100f8aefe20f40e2fd4f71deccc",
      x"6fdd3f4eb2fec3e30a04c7a1ca6aee400b9137d863a9abf94a7efca74fe2cb62",
      x"191170fa48b7df3ab6c19927b37df8037f9aa7710e8a727711077431c70aea58",
      x"ac895e797141dab258bc3145a320a4aed2ff136a57e57420fd6e9a4206f9a0db",
      x"82752b5ec0eb33576e98a1c30d4dd55d38190c8b8b608570b632b1173df30f75",
      x"6382668ee5b94a7e042d0703cba82dc5c3269fc957046308ba0b7cace2cdcd21",
      x"05f4cee06eba13e3e52cca3c288e73e51ae8c7a4d2c731319d9aab5c8f679ce9",
      x"1f4ecc6e49a674dcf02ffbacc5e35034cef27cae3fce1f297b930b30faf82cb1",
      x"0f874cb624ef0ce2a6b31534c06e8da8a5603c8947a056c70d419e85b82d7f31",
      x"e03161f53216deddf7876273483a62409a975b8c85153113fd7dfe0eb8263237",
      x"e4e2352680b71e52ffd19987f25fb33701239932b2706317afe94a93483dd79f",
      x"09a9d9135a2c5a8c0c09080a77971d7281fe6e3f5252dceac87bac897e208346",
      x"b3944b3a900175fe05dd32be4025070cf73d21d1aa5e2b15be37c0b67fbb0186",
      x"11529a00db0869859e239eea265dbe4e049d2d9e0824927c379ff98dfdd35bf8",
      x"c91e45b908d60bed6f9799f7a68470d26d6c2bdf78acba729e94310c8b08c06d",
      x"c5e5b8dbcb26888bd8eeab94410d5183cd1b70df6eedd076b1eb789cee97f187",
      x"c6d1b565dd66969708537075b6fe0b6e6c137a4518e4ec9a495a82721339b41b",
      x"78e6c87b97923f99f08d98cd864885a672f073214a1240d5f856fbc0b48426ff",
      x"400d70f01c81120a45dbff5a191b26bc9ac35be4480d278b3e6344c092b7bc11",
      x"fa320d4a910bc4b0d7b777f24c6d775bf930805bb592d8278b333faa763c7dda",
      x"6ac2711ac147df21ddff588d78b4ffb781c3521b2d18049bb744aa3b2244442b",
      x"c4517d667a782e0b9b1a8be96a69458d801fa37d865d6a579093d99224080ce5",
      x"b416f74ca49a98279ded67d2131540eebeabc8c6dd39208224a1226cfbb471c0",
      x"bb12d62cb8bf70e7b6307c89ab1669eacf4fac95223214bfc4afaab72c1bc599",
      x"66988d441bf3fd793bb30d0ba60d4e0637b2d23b6631efbf93d8293d36f45e63",
      x"babb88a1ae7fbeac683b09cfc55c7a8d87dc9c7f5d27e52af82412a9a025da84",
      x"96c8c8e806954ab746a41d2e81ad37b81f3720865d169c7107e24169a20eac6d",
      x"7e449d2a4a7ae5bb0a50c406ed521435a763c7d1ee4978d8eabf3858c9ed7a72",
      x"d2bfde4459e70e87196da7c009cddf4b04f07ee06044109e55f9323dfcd5d545",
      x"e75ef2c19afcc75d792bd3cb1b6f56efff5591102760e27aee4f2fd285cf08f6",
      x"44d75a243402c845f0b47bcbd8e48cc064ad8437c9d79ba0bade92121805dfaf",
      x"2a9ff53506598af384d2136f392ecfcb83297e53d0731eec9b8143983c4821d3",
      x"cd71ef342fb5d8d0a39a5ee3c6ddf8a8939ec2438a8d4e36a79e5efd31a1edb8",
      x"a3153717b3314b2ed5c9141227bdb7ba082541fb7ce9d5557a07443dc420e4e6",
      x"45dec119ba0ede476976a1a4154bba309b755425a225ddf7022bf1fb1d2fded3",
      x"b97b91cc3a9328fa4afc36562d9a53931d084c8e5561354cd744d8e7f9c5ce14",
      x"25ed3a0b7c46bad4fd7eb050971f8ac45b49487d5ed804b98b8727459d21fd11",
      x"aa15b64b4a7f836c27a9b1e0dc10494391963963b2b7aa9719759d1b31b2112f",
      x"3b4415265962c3fd0490cdb76977c34037103b16381837afb90f455a017f224a",
      x"d2a8eedab6242f7db8c670accdfd7b195287da7efc3dd12275f787299a5ba210",
      x"0917373a5e1911f16d42b3b6094de9d63eebcd3d48852fc89aa1d882a8f0d00e",
      x"5788b851f43694109ddf95845cc907e4d363cec8ef36a2718b7c7058c88f061a",
      x"b95177e9e7a19ca74d18c7da73df71e2e97a6862aeeee30533937c88b2f63fb6",
      x"194dac560f8fceeafa01ed5e1d3c44f84307979c2ad2de2fd3b3869c8538f43c",
      x"15bd66e01900101388cf30ee4725ffe2e85d993125f35e426c38317b848adec7",
      x"7da0e380422d13b0b25f3b5ce6bfca04c6e1304f9f92ff06314a50ab3eed06f2",
      x"e12bb8fa5fb3d446db8d8131ddfcae3e5274220534191f7d046a0b31e055d128",
      x"9a74c976e63c9afeaff4488ac940621e35cff7cb3f0d4bbfd5bc20e741a8d23f",
      x"62658a574fa444f0762bcb0a742833eb7700504dda5d044e8540e74d796944b3",
      x"e58d18eb49b9d3a8d740dcc7adeb70777182ef5def4942421bb62433e7c24af3",
      x"6207ab78338a6d039e5479529527f7b13ad6463b0f02044c4de3d85ad1ff1e91",
      x"6ed6cffec73766cd50e0305af207aa5137ccd1163d45a5d2d18e96bea9f22aea",
      x"d75dad19edf8477d4c709d169a964c308714880af81b413f145041aab957775f",
      x"7d5a13f67fadb4489416f0c3ed80b97823df30676640500abc1f172485e75f20",
      x"005d153baf310400b295cb2a2f1e1d7b7390e762554c1a392fc4fdbf8211bccd",
      x"c9c98c2353f9d8807c7710b90485aa24650c07d084067b93b60ca6e9c7a4dbd3",
      x"b94930157b6eb0d9b4b40576ed08e8e1d7591c431937af53211a024cba9c12b7",
      x"b3bbb813726241497432810c8a71eb436563478266aca09a8124e251484ba004",
      x"be7433d5aaa5d224557ea30835443f87439803e420a1cde871c97dd0e7518035",
      x"6f9feeaaee2b6ac67b412987b36719fee5415d21ff7d82f932b55228006577f8",
      x"3ca088ac23fa2a88c57cd46a38afc8798e147906fca7ebfd650bfcad465f8380",
      x"7e149aa6d1e6492bac318c57528a7128c7a5ef34fec9e3dac27bb5c43b66bae1",
      x"ed09abf13b025082d70336f3faad139d478b62f6bb7883e1ede0c743050861c4",
      x"9ea8cc511a1e777a78acf6f764f39ea2bf549594dce4cbd3fad090df7f2e1a2a",
      x"4d4e1dd78cb5ec7d80abc8cfe9eac20943e88c80b5baf9439acc584371d95d1d",
      x"187ce88ad982436044cdc456bfdddd9733f765f1507bbfe5141ac6f5674391b0",
      x"2926170a1083cbdebab492ea01d21282dec37ce7a3b8fde1f48af1d51be74806",
      x"ee87d091e4faae70f39d66c848abeb1101c72f96f972809399f492f11814796f",
      x"dcd89671498fa1eca01df2ff158a8ad547fa8dc92497d6d94bf6c433ff808a14",
      x"83cea3d5224fe685391d1bd809282fe159348b59a9f49184bf690faeea1f0e04",
      x"a12a5a476b1125f858448bbd1b59159c93254105501850533e3362d6f1738567",
      x"82ce9913f1382efb6810bd345a4a419abe06db836fa8eb1079d3c3566a3a7493",
      x"cf8c4345672d0f0e1ff8e1b2af93cd1cae13a98f93703bb3644dc63c9d4c8493",
      x"a5926a29bdbdb784bf51fa5c866ce35042c74dc6c0a2e6a21500b8e50e21d115",
      x"1d106c4e18d2ac7cc7e1e361a703267515efedf549c23eecb413a0b0847d5eb8",
      x"4f188de4fb82fed9bba05d4079821fa05bd7076f3e50149f523a73fec4ef9311",
      x"51b9ae02d916b847e8336b9ff2849e00fdf9ec0d379d0ba588d0c41afe46a8ea",
      x"1ba8c252f2ed679e73663582e6bed0b4ccf34c116af4e49471411886407ca370",
      x"3b02ec5009a3579b6beceac632e8b45137a6c8616da274fd9bd8ca911564a708",
      x"8df5f463205720863e6f865e09ec3d3e95e419b28b190913923d12f00f901710",
      x"37e3963d7c1eeb3c3d8f496cf27fa3833fc7a6217d6fcd16de3e39ce4bcc0024",
      x"dc9e6fcc1561d62d22b77ba40c9256a56281b1739a271b5ffcb343029b7ba388",
      x"6bf3f24844213d6f5486d51bd384e1652170ea0f49fb633de2cd2cd420112638"
    ),
    (
      x"3ae0790236bffe03a0c5ee08b583efeb76b83258959262c29b72c2056756c12f",
      x"285d582076775bc0cb08a30fa3ecb0e360063cdb47e50555d46ab797cb3b79d7",
      x"6a2546dd5c008411dc7a565230c201ba32e9d0d0f53ba3d2b20e2291dffb55b3",
      x"a4112527e7746d2b8f954c8a1adba1e33dbd0ac0057a2870aaac2c65a45d616b",
      x"7a40488fe0f49c1c826a4a39bfeb63e9e7e5ed0bb975866e8f24a2d6c47a704d",
      x"1343b8525e5dc417952560c455b52fbe7d3d6cd8d13d76ce18eb5be24c589b9b",
      x"81b9258566ce97c961cb53b54f3f14c1936074249db86fa64fd2e663a67489f7",
      x"b0f6b861fc950e5fbeb51a2f93d34f7fa2eed2d58b1048a55143e57b0b840e85",
      x"ce4d01b0e4b5ea6d27be2801661ab1168fb6051248e51e8d8e0d04eaaf86227c",
      x"7c46bbf57998f5c28754602d2eca7392133016c04012a54740aaaf4655c540f8",
      x"ee420ac98469fc3c8a3bc0a852b3a6a0f9e5753759294904eedd1e126080b9fd",
      x"24e6c02874af2bdacbfcf4abea8b3a7cb8757f655f1658cf1fde5bdffe65e5e3",
      x"f04b55e2709ae5e580a802674ca0187398b5d703ddf9c3352a43355a7ccd7c50",
      x"c7863efec135328b18a740c6662ca882f58faac9c622f5b5b5c8ca0bd0aa5a9b",
      x"d1d0f13eea724d98b791347ed82eade7c1013142d8bea0dfcced637c0ab8175a",
      x"924c575dea3ceb069604f65c094c52eec889c0fcf7e935405a31c9c47ef61766",
      x"365cdbbd0b2f1256ef2f4bfa2854db0621f700be813493cb026a78b1428844fe",
      x"65e3b79a4585e1b80eefd1d7354544497f3839b57047ae4917f3cb41206cf5f9",
      x"04a61e238d72a09f5045284796b021b0a9741a34e2a22ec1acae322baf630a8b",
      x"6fea92803e21e820bcb43cd99696ef9bdc36942e97e522a75ed195850a10acf1",
      x"694c8a04b89fbf237a6a8c528e99aaf024001c68cca4b187a459bc859ce68e3c",
      x"d392fc76046dc857f1f355dc776f7e18de27a2be78fb6112f0d8b6b44ed80914",
      x"565b10d3c4b7a6a33e76cac1faba6139eaaa26936147b9723c9c649d674fc9c5",
      x"0571958999dc57362c0ea46dc5d08febbd6371ad89ce3cf5fc5664ce5d924185",
      x"a2da87fa4c70d602a7066a34042f83fc0c3e8d079459df0d69179e6c49462371",
      x"5053c26483eb02e8d0ce643ee3f95bde92b378d56d3810e4422ada042b817c6c",
      x"afda51ed22316ce64949a6c4c90bb94d2915c0e168dd6bb92c0eb11dd6d0486f",
      x"f162cb17d78de960fd2c4c5eed99c15084b9ce8016425a568f74513bea39f872",
      x"aed0c80641b5588c7cc48ddcd27e0d09a8e43239c33d669f43143409087beb98",
      x"e913ae75b388388dfe1edc1d71bfcb78416124bccfca4c58e0f8be26a69d5b7d",
      x"f04f73924fb7f8bcd8bf844238fd93e77395463f8f64c8a3d508a6e61444af63",
      x"d4913803bb76816d732ea02f098c04a46326b3d2ae72eb1d22b2bf73bce315d6",
      x"2b1518b06fba0ca2928dc7585cd3addfdf5b645d2461be4cc773a27f39d15a2d",
      x"99aa742ca966b6df823fe544c5ace37979a3d92cf821dc50687d8d7cab35e00c",
      x"99b4fa956040212122549a56bbe78d7a7051e60c34450de9385f6ce50f109bc5",
      x"1566fcd4f75b59ab4306c70bef4636d823ad71caa3d3ae391f42455cbde2fc29",
      x"369642156b590f9f788c4b639f20a59f5705fd640f4f1f3c93f9a7450f2a5ec3",
      x"33a25de7d8c48534ce17d607e1a27a34ee5892389531a844e6bcf3c17c22e895",
      x"2dcc6b18e8f249163735e7365c7ad87a320c69a3849a3059541b64c88ac60100",
      x"0d82823eb7244d8dce7b31301283d4869cde453d067cf9faf8bacf025c9c6ce0",
      x"5da56aebd657e67f14ff5a2467fdfccfe6bfa03f4fa3ce3c793947672303b105",
      x"f2b85cef0a7bef87fca9f1f39a8b820d613ff67d8e30b12469f50447b377309d",
      x"ad51161f37f1fdac99e67a72e22bbbaba39a9ea61994fe843a3713e4ae803902",
      x"d80cb277673786e98b79f5c8db0eda23336667edc27072bc4aa9c44dc0a1c71d",
      x"c2700e20d85f47c20c01b5dd2a6683749ceba75f0b4f6a9167885f31a6cffb49",
      x"4719b85f4c0aeb73e37e5a6727def1e9025699824eddeaef2cd0dcf2616b1ec7",
      x"0aa4e18a165b8821103fd73a2e3e7d93e27a920cd4102faac4fe042bebfcaabf",
      x"e39cde5693c470dc4c3e15b144bbc92e6e6c726031a69526ea2f14d2dd61c845",
      x"f4125447f352b272e97e88f957d492bfcee7ce9d52e2872bc20bfbb2632e0e8a",
      x"cbde3682bf108ab97a4b7ff5a96f43513e2fecafc1f4fc31bb051e14f72b66b6",
      x"49ac8e6a9ade776cae383cff5a3f76e753133fa2327e3bd52d3d95727db6efcd",
      x"0e7e694a5075a20421cd95a974b5f5e3f1905eb43808ecaebced0989e641dbbe",
      x"f58fd4d56abfe2809bcf2d2c1fa9605efe9b8d765a7baca042c2a63973e5c71a",
      x"c429952445495457e525da0b6b6fa45dfff6dee1f46b8960e37ec85e3f19fd38",
      x"293238ea2c6321443e2b875c9e09ab221ae033471cb5cf760a3658a4c980bb1e",
      x"35ae25f9192709b06caedb6280f7dc58789fa9bde40767548c5ce9919ea3bc6d",
      x"f06c233a431ebd1addf6973e8130eca39bc5a9ec419e4dbe53fa677cd0ba77fe",
      x"1200369a6216607e4ae6f03bc60712b0468a45aeaa7773c9fe0fef1c0d2a314d",
      x"d6c89102897e876cdeedc1a1958f87c0c3b55f0401cfcde8b11aa32d33b2f46c",
      x"e92e316e9d9a47b0f07cd55fe93f83ca9a97a226c9f3a958c3ee8b509451531e",
      x"fd6bdc23c3874ec7233da94a8a18e0e24b199821c35837881ffa565747dc02d8",
      x"76b7d2773affad09f26a5df7d792dedfefc3dc9d81bb61695047b53d543dbe74",
      x"572e1da8c707b71a757d67afbf84dc88b16219acfdb1a1ee867956e04ea44f71",
      x"23095fb52a42224aaf3455d883951cc3dd9aea52a8ed2f54d3bbaf8fbb4fc729",
      x"97387d182690af276832855ca241bf6f3759f1e0fc5e6d18a3b09d2d4f096b9a",
      x"3d1b2070db6437ac69fc1f7f0ef3b648f1aed12551a53ab89d0e0c3a435ae20c",
      x"52f8fcd2267fe927a7cd5ff72638fb7c72863ac49d1809cdd408accf921523a4",
      x"40677e9cf888cbede63617e1cf1b68938f6fb776647dfa693e200d91704be9d0",
      x"9be6c0492858a6cd2e5ad03b606191d37f58f2ca448fdd3b7e50d1b20225372a",
      x"6592a875e4c1f75fa8ea69259093bba3413c6ba7952e33dfeae6f14cb6d5d0cc",
      x"49299b9f6d1d3d750db3b6e1721aa084fbc1f49c1531385007c3e3e60761f843",
      x"91e6a49df477cf01b8a9d0590e08ca52307dfd12a9ceec3904491cf636f0bbcb",
      x"e7c0cc8bc2ccc5540d8fb6f8a2c20a4f565673b8ebc19259e7dfc68ff084dd0e",
      x"dd6eee72849a23a91d1432063e67b08633eca679de2ecb5c53424ef01b3bdd22",
      x"2f0404de4a76bc16662e47981a54aa5ea0ba5ec6e6d6609f2726c0ed9eebc059",
      x"41ec4c2f0f19fc6b3159417faaaa17f9ad5a000f72a717bf64caeb1878628a36",
      x"68d496111f6ef54cfaab7e93e5933e8703691bfcf5e5c0c2f27ca24423ec1822",
      x"a32a1d34fff3b91d38dbd4376b05af11f0b98862dd53df0cde3786e146b01bb2",
      x"a369ee331cb97ade3f25bb398ef9116a6b8d47371e5af58f6ec6b9aa9e561ccf",
      x"4b48342c6f5034f8a3e9341f9382dab9b6677c0fd8aba1c484490f18548aed64",
      x"a46da7e78ca2ca188ec6f7e8b1d78fd086741de30968165a868f499d88d7db17",
      x"f194bc2d73b1932f71bd6523bb8e083ea5fa50add3ae7111add0c25f79fd9713",
      x"a9c30727e06b73b019a1f65e07bf5c82b3938f0b7df9f67e1e056bdc3ca8c1a0",
      x"d88fd20c27d3290e6a0b113df6734b0b3057edb878613f459690dc2df3bfdd68",
      x"aee5302353d05d9c2d87edf4c9a3b94c4b77c60dd146822a094db2ea1d8c422e",
      x"c37a918c2d69ee12a99cff0f5e2558087a202ae69a526d36976d985d470ba34e",
      x"c0b71bb0b4f7df03bdb8469db27c48f09e6c2250b9e7c4d6f867ab4ebec7d8fe",
      x"8e591e33789d4e9888b6b6e69fbd78bafe10c054ef1650dc305306f587ac0ee9",
      x"296b9b9356d55318c483113b6f0455901800c04a0f66ffde690b668d0aaecd43",
      x"06678604edcb5531f96534794521b822d019085f9edeb8d6ed3960db9e12c93f",
      x"7b180b812d0ca67415c87a6bf169cb2fcb738196b66d6b5d58fb02667a2e3a08",
      x"c74067ab2a301022e4d29e4b06528da136fdbd927cd9a5edee68dc8231be8e33",
      x"5580e286cc4f0f73d9212a4c3233cbf35921e322c4f7713a1ef5b919b6a24504",
      x"b36f350429b9dd679e89856a8bc871ba8eff02aa37df16927f229f35571807ba",
      x"decdaec45aab7c79692f75e65d4c460972a64cce7e6f121640a3c7f2d1d4e752",
      x"ef5ed7505a192ad4780d04ebba55806cf3a6ae13645e51a810deb3922a7dcbc0",
      x"9f2462b6582be00f25d83dbe14b3feb624c7f92bc3f1ee2e02f1a63b6de0e2af",
      x"ef949c4dba49dfa179ac103bd2834383de96e68e266f8372c59d192872c5607e",
      x"54a273d3217e25c4c01cc488d8e11878a4a27be99e81394de8647eabd6893a88",
      x"0de8e17f91690157b6ebf7b084dbe8e690f04ce91c9abd14fb1589f248023ac4",
      x"9c5c852f4a32d1ec127edce318266f9f2565aaca3e3fba57bb6a1ba262a983d8",
      x"80ff18dbc9f64d94d5e616890990d66be9d3ab5c1ef6ef0eda091a9b212d74b9",
      x"dd6c2551f6bb0f9fce561c47e2821552a278224a63ad9f380e39043d33ac891f",
      x"789fb59069c205e12d2f9df87863a5e151446c86576d0762d534e080b7364fb2",
      x"739475a8f7a0ff0b5064f50b70a8bfc05eda2dfb8b123aaccb0b95f7ee28047d",
      x"26094daedd714ce3a7007231b64aa099cf6c57b363d01fdf5bfe4cd995a98017",
      x"34e6e253fa4b87c9a1da4179d997b91d322985d08f81a6f9f4943c7035a80b3c",
      x"a8707b3aac910697834ba12f8ae6dac61258eb5bb17457337eddd34d26ca11f4",
      x"7894e9091915863494be510f0f3cb009159c64380c057308d6b5d6672e997731",
      x"442d30dbfbfe14d6f4ac22472c84f9fcf45df2761fa72c8861ba46794a39717a",
      x"f4c958b282d7d89aac2e93c82036a3799175183dc0ddefbe0f7545ffd84fe2aa",
      x"532842d3cc4afa3fc3ca4dd0a33504ec59acf0351c0494a29842861c9348ef1c",
      x"6f159470d0ddef0510861993a35cd73898a149c6df6b065cd37da76e29309288",
      x"74e7b31584cfb621778a0870d0c5d3de7020ed1ee7036697552a20c263a509c4",
      x"45ee04b60c5addd1a9ee701d7ca2ca00d9df05f682ef7f0562186f7514ac4ae7",
      x"8844a3b7b54bc93aa217287a47d02f678e320c08fc9c96f3f8fc0cc0067f56d8",
      x"7748ebc68c1e5b44e728dd9400d9d824f3341e28911e5edd00979b29d25af5ab",
      x"b09fd116db2457e3c72f8e15c9bc68f0b287c78d640a2e23f564ec5ed99d08e3",
      x"2c5fd33c6a42dea17b848aa4328e95fbc6731fc52fc3889346d37d395235a816",
      x"c44117896b346ee4622c863ead8d8854f2340896331974dfda4742d66635104a",
      x"c9ed63584778e956bda1594446510393f9082292ae5a9d554313fdee4fa24b67",
      x"e8a64a2c6c4d7fc71b62dc4e40e5ae0ec5d36d2ea67a8a2346a1e696abf5bfd4",
      x"7c2f5ceded2b92f82f016ec0518cba2b3207e1065a000f00c9e0ce2fe9b94fbe",
      x"30053d967b5f0de5d7ff4ccdbc9545759f257eb5699deee4c744ce3901aba21d",
      x"be1ce2b858400b2064c4f27cf9b0273c291ab8e242eeba46412dca721870ccda",
      x"519eda12dd19175576a94dbd81ad20cbfcbfcfb32cd9816d95e2aec035f95fe4",
      x"601f92dba670242d0a1d80f04e24d53dbf12be4d4e2ae0161892657cc9d81c2d",
      x"7f0f40068f745b11f941bffc3e1731e909f9d9c868318fafd017b0578e74306e",
      x"b7fc046d5f0ad4ef4dfd1388b75c2fb81b05173693e004383385c3b75d79418d",
      x"4aec8e31e486c1bdaa336253cba9ed553aa0bffb298b741c7b632bf8014ea12c",
      x"1c80e58ea368db1dbbbb8a448404dbc5adf8a4b2e3bd603f756aa157ce8b16c7",
      x"5a70c9d0d25ec4d8356976df072fb24158ada6a0399ba09d1d90cf10e70c6f54",
      x"367111c089b14d28a79dc5b5a10204ae868da85a3b42e1b001bd8963b42d8f2d",
      x"d1edcf7eb1e9dcc392e28ecc62b762029d8fd68df924034334b069076a4acb62",
      x"71385ccfcc904dd9006624020e028f9b4c50d71b7effbbb280dde8de742cf8d2",
      x"4c21564ac265976fa9631ba42b7205a38027802787b30a41f6f4f403d5c82027",
      x"7c646e5e197944add5e89f04128fa70e02e1b0212e64abba7fdf86d6fd94d624",
      x"f016706ab1f9415e278158718987f3ad466b458b6be89fce28fbb9132e9cbe01",
      x"0890982784d3780b79c6fca55810a13a4a9c42435a4ae9064f59584ab535fe85",
      x"4b7116f0a8775379d2f535d071023d7cf406cb951ac6879e66a950d6d8fc136d",
      x"7edeb393040ef537c03183a5c6f9c5934c47ffd6be503dff0cd832495389ffa5",
      x"45cc14004ccbabdfb8a6c10f68ca644fc1b8336086f32bff6801d42df5090a33",
      x"a3f04699659b41f093ddba664f746f53f11a74b697a17fc97ffa78439b09f1c7",
      x"9252b03afc4f244284e256daf0ede58d2d0ac9294840458b054eab627c8c8971",
      x"8e89e2455e07cb1714577c6286392fd5560b2d0f7b1f1506d716a6b000a5d058",
      x"924a100aa7bed816c3b939258054a1af32ed3dcab80b6a54add96fb0a8188734",
      x"c6b9e3d2ba626e618a81441d0fa05e6b9fb078152939763241b74cd7a550308b",
      x"d729308b45f3ef81ec0a8fca0d2f79227127ed9b65d592a6579d24ca0b6ea405",
      x"0af1fa0c61e3eb113fdebf4656074be70cd3ce82598e365db6e6afb4dd262160",
      x"3f49089543a38c93389055170a4d044f30a4ebce531e6c33aa7b123705dde2b1",
      x"cb3fc57f571a0ed08c0b3da74dc5afab154c7a3556d8f8fee3c17d9d6acb35f0",
      x"43bbe11c70a656ce4f0f2b6b4df9364f7e96a870279e0f111b2b0fef8b9dafee",
      x"5d8b9e5547caa3780a1c1e122e0f53193c5cb593e57f4138d05df22cd3731d82",
      x"f7a8ae890fabb3966dca0f46816834993ba658a3fda2f9ad6ee00794e313e9d1",
      x"901bfafafc791809a82d00759e5750e28f3e3de60354b9fdeffaf8ffeb875b11",
      x"4900b48a63d6bede6999b8582559a372e9baed6b9bdf0116085ac0338b6207f0",
      x"8a72c0e23efcd076103f44cf7d8c5c03a4ab0f7c7fe5a59593f4f9e68f37daf3",
      x"bff66458eeece5f6be5ac13c36f11d9809cf674c28f49cbbf31d1cf7fbb5e792",
      x"dd57f498c2d1714315d578913a8a948ffc42ef32c6cf2e9802dc58dde568f7c6",
      x"9307721c3d66811a1e16ec84623fd37a209d6b9feaf5495ee76fd333d35b1d92",
      x"4d00cb1b92964e8313929e8c9a0e5ad805d06169cf5609f3c26e0fa36b8590d8",
      x"118eb832f0a8405d0020d6defab7d35db2d157bce2c904c9c8201d3e98a8551d",
      x"f33d8d17d119fdcaf14c25dfe5c147888ab803c5ad05e7e61a0e29c498a35a61",
      x"316d0bdb982e7b8a30933c5403161b2e44a907fa62279f4db38b91d67bd23f07",
      x"7792b29bd0298c73519bb479221e600cbaa2ec87237b87c945ecc3d7abd8c480",
      x"a179e54c16bc545932ac2fc0a9546651d6222ed16034273f124043f3a11730cf",
      x"a9a3503508445f956ce8df0822452b2f9b829d552add592b5ff16e789f0e0994",
      x"7c2eb593ec8818bcbaf39a2f03b12c18e6ebf1835c782eb85da5de0505b59f66",
      x"547e5a1f244752ed7861128100629d194bfb9a58917f6c339aa920fe4fb39a0b",
      x"9e9cf33d0019b2c5505284085463fe5ed135ffd3ad35cb673a021a6837f6c3fc",
      x"43e327b7c4db48bf4bfdea26d0f050758e92c5c1da09cd2ce34b4bf6e6dc0859",
      x"01008977bf519ebdc7be30335cbf9070d4377a68b5d31bce29cf50335cbf3c16",
      x"08ed68fb1846b0a35db096a54b25fa6fb54f9c08d6ed86f6c58cb013c602ca15",
      x"f0e6738dd3ee5300b347c75be4fd5608b6573ed4caffb0fc2c52ce5610871daa",
      x"48713a2eaf1cb75b56531d426a153fad943d365e65c1c223d670b000e18a8979",
      x"7f21c32a7aff6130c35bcd88d1293622e54704753244ce3f9e8f318447d13af8",
      x"a5a17315c405aef7ee9fa42d1f536b07f7727110a449fb47071bf2655c2f2272",
      x"212b8c89d94eab7112dde15f74f99024d07bad83868c54af52dc4945de8eb31f",
      x"504be337454451b111ff14f9d25bfc717c5b9581204acaf89fa2335074b1bca2",
      x"5c50f8fa6c3d9cf1489f00183f40b1d7add6d4f0a1f11a9a509d2eb6f94f0c65",
      x"05ccef4084f3ff501fa17d6a1bbaed1fdeb7cceaedcf7923d1137789bc5926ce",
      x"0c808666deeb571704c4816d74996ac37278e5ca479349af6256764646221d78",
      x"1a9d5cbc7d777625a43724b4939997b8ae0db5d8dae7d4ac0ec90097813a6547",
      x"cb7fc3a5b295551f5140ba8c8b16eb093395b3c7f093cfa2ee89104966fe254e",
      x"6b2675d51f68d736ea491c55f9dc27a6c6ac59a35f847db7630b1e1c5873ce40",
      x"971de625d1d9d4689e7c9fa6b90acfdd9283390ae5fb1e1732355d3ab29ce0d4",
      x"9fe0e286c2ededc6796717e0710c607ca69500079ef19ffc00ee1b0bfcea13bf",
      x"7450f3493b0ea4bb30612be6f92eb1b4a757202e864deb0afead19e9057c6d48",
      x"4a44174369eb5cf1c070fd06da8c29caa563d3dd9e185ddc9eed749d2e2dc99c",
      x"653d333839fe0178b1e08d59618bcfffecea8f8a5dbbd1295929080d4b1bb09a",
      x"fa8bb6f8862dc9a3669de0bc674ca32e81e2475b40c43261f0a10eb8e6cb2438",
      x"2850d26a385f17246165aa5450e3339139ed9ab4578fe9c062bf4711940b3036",
      x"55f94969c4b1d8d5956d3a5209fd7d53ef3ea100c58bfde9f83a2e12c5fe417c",
      x"518da3cafa0dda7fb5bb939460962355fb80baf03267108a2f4d7c55fd19829b",
      x"d17007d87250d0ea670894f8705cd9d33ad43db3ace6d02bb75cc43f9128d858",
      x"12f6ef0173ed67590fe94543c469024c8bdd95cbb045ed6977e05f6d45de56e9",
      x"d594369ac30757398c7a72cdec785b295544a98875fcee859459f72e3df57ccf",
      x"a3fa861c76c25436236e1781cc798608ace9d2d2450cd47749c7bdaabd623412",
      x"cfe0badb6bff89e3add312d201dfec3294de86187d15716cce42dab2d10bf3b0",
      x"eeb2966755ae2d41b35a8b139a5c9dfac7e83c0915fa202ced0a70dcf92ac3d1",
      x"8a746356b7ad38b77a75995dbad0c2ec2fc5513face4b5fc43ff2b0b75a3a38c",
      x"2f47b943fd34d3fb3780b62a90527baf855e9d9429e71ae4477be583a1dac444",
      x"a8d764b08c8da399b9c0c0b2fd8870a97b2d2b39e4bde53df953e25e5d2a1f61",
      x"538e390a9ae338031a7ec49824e888920d16f3d492817f5fcebf7e181da1e27e",
      x"175816235ea3b42ddd186dd8721bf2f714aa27bccdfedcc3ae45a1cb5dd565bc",
      x"a472351584e4dea2267338f0d7602b15cab937dc2129f6cf4614ddc78dc7502f",
      x"053f8ab7be530b878ee1ce3303e9690780c55d83160f0b45307f9cc302b8b4b1",
      x"1b60c3256732117ea2e74421aff10f269b7397eb642790c4f0a06eff55fcfd71",
      x"bbc4fde0e798c427cfbea099464792509fdf725cfde7175fda21c036d81622ce",
      x"583160694e1acfa5757f29db4137726ea351ceda6582cc39b89cf795a9aa160a",
      x"76e1ce920aca671fd3a74ef83a641dc7371449fae6ba159b8675c5ca6a65fd07",
      x"e490a5503b5eae113d5f98f8f6671e6238ee94b1cafce2a663a6e64408bb1011",
      x"8c1a76f2042e1f8fd15799861d328fd1393e77cd051782e7430e070b4f9fa134",
      x"4dac206bcfe53f04caa66793e905b7f2299cfcd7602b491aeaa1954ed034e82d",
      x"297a0dbc3f176cf26f873e17f245cc7288f116648adf8c0069a2056b49aba173",
      x"1688e47e64ccb2878d99c9b0ae77303711cabbc061b67e5c3f450ceda2a81994",
      x"b5faafa105d7fe35680dc80140e163b63cbcfcb0d5223f37f7a413567790d4ce",
      x"4a488b6c7dc11d13acbc762fb3bd059cef376b01aa4b63b76941418ad543fa7d",
      x"5a2e3f6c2937a2522f5a9ba7d7a23adcdeea9d8364a827bb398b2c29c28f11a1",
      x"5019538033afeb71b76dc94d7ccddef4a17fa3545d19671ea13b5a58acfc5145",
      x"52665cead1189fedad621d24a185df69cd48e8e70bf18b1f6a874b3ac6bfa100",
      x"8d187d7c2a2d275848b81fe40b2ba5b01c19801113693b921f3fe9c43b4339fc",
      x"0ef2336f3bc547ad346cb7cf965b1eb8772a3e9e554169f732cb64271ea7f1de",
      x"56264751c20dcc4eb105863d1d42feafaeffd0a08d14ad6d0ec19deb1e6b053d",
      x"84223cc548ea12e943c732672f86d8d06c22172d7791ae297c25cfc6c7c29272",
      x"92d02307178528b5749ce3f2aa64f14eeae76b45ba14869653de2a42ccb9d6dd",
      x"4a2eaad04dfd7db12d8a672e2d696c69847d609756cd789f90f428d3e744b711",
      x"4bc4cc5625b82dfa98bb4f60c70b0b78c003122af66b68bf1a2f182458e7aeb0",
      x"9ca0241ee134496364eb3d596c25936736e1a7c9965217b8c56dcc600c6225de",
      x"60833b7ded8eb5f71bdd9ccd474460a092eea4ecc1a56c880b18902244bb2afc",
      x"b148d5a667954036e85d8a74ebdb1bc076e25009c2b50a6bb621fbec340a2721",
      x"e5407c9f732659e8735e0a97f01953f352a44f92778b3f7579a45d2ec63683fd",
      x"40f1a84027f4692a4ecffe305afd224f852efa3cb50616166976ee6f2f8dab6c",
      x"a3e0c714c66f815b4bdf7bc8ab9e46442d50abeb2319d4dae01eb884e8f328f6",
      x"4c598c8399c8c39498f94203f0cd37e22e532a98241a99214b06f4b8701c5cc7",
      x"73abf44cec755464df3409b268d348a8e482ebb902b70b56de65fa866bfbe609",
      x"056d26d37057ccc6bdcbba13f94528144c3234529a552845e54ed62fe7c32293",
      x"fb3a7c40574484666289fc975088d175668c906a2bda9015f8f50d76d7caa9bd",
      x"9ebab9fb208f16a31f7654df9aaf170bdd3cd4d2131ec12ff77511421670f60b",
      x"695e454a35c5de655a7d7e71df1297a85b6d6f3b3ab992a884573e9b0f4b810e",
      x"69545ce582110247930bc6f7f4621ae3c9907089ebb7cf4594850c510b155614",
      x"170e97f1858766356c02b7a96e2605d0a58f06409f01cc296eca1620ef23201f",
      x"15f63cd8ec271d75072a504eb7b3bbccb306577c2138749d827376341c88c36f",
      x"a4901dc15c60a33684660bc672d85b3ee996d9a6e20395c6ed7585e600fa209f",
      x"00ef7e057337931af4144c4dee44ca96ad913ec0678a014a90f7a8ecdf3f6935",
      x"415e7b90436e0d073a0da954561261748681a87748f1e33f10720455633bc8ac",
      x"7d12eeffe6e4b2c4f11643faf7227450a013c0bc64a1f5337abacf106d8ce9de",
      x"230dc3eb861ff67626247fd32ec613ae4c6dbcf781e2f9008bb9a76ec845f71f",
      x"36a33272dcc10732f3c8f035f13fac4e15fa39d390b0b7fa66ddb2f121afc5a8",
      x"0d53287694f9dcb64c347b5f1ce78cb821a7a07748c61354b68a832add990d17",
      x"9172875ae2ab20fd5080cde3e54814360bf807defcca8276d41176237a76a505",
      x"bc4155f0ae5bbaf81c01ab3b294ffa02678ea8fd9fb95ab67e023286cd53539b",
      x"e10d9c8e92f33429cf9e0ff8b744fb351a06f95f78f63267bdfe05e18509e383",
      x"d6197226b96976375ec453477349c5dc32a4c3f2d326260f8cabf3db9af3e29a",
      x"1675564914eb99e10d46e22300ba0f9f0b506da388fed4b3a78ca35faa6006ae",
      x"f9e47575603328da3abc4a0e0487facbc4981e75a2fe8597c06c23135f195f94"
    ),
    (
      x"afda8e92f5419923ab3eab5cc50fa7f080ebb0245cc548026bbf6c3895860275",
      x"034aa964fd7442d2a12956c0aa947cb28f3e3cd6d34c2d560b8a4261d8b7ff9f",
      x"84818effd6e66a97536902ed33b4fad9baafed1a0ee108f4f74be097fc16b8ab",
      x"50b57ce0e55082b52c8c2afc8f4789fcc423b194fc586ac339421a554cff4b99",
      x"0bf123c6d21ece404a053a1d7767d2944eda84588e138e7dbaab44572bf3e990",
      x"cb14f08d53e40de7e9ba412700004aabe6767cdc70e76e0a3f79603a18b737a7",
      x"d7c2dd10ce59706b21222854115adb46bad82acb8d91d4fd2c6a1b888b69d709",
      x"ce73248b6aeef0a8487432b9baa9d1ffe9b2bb47d5d6b42ed02d1efbd8e74cbd",
      x"bc1a4c09099e2794cd31d92e62c6981f43262dc58cbe4d4f199c1f3bc27a9834",
      x"fd9205ba7219a756d11a8bf95c2681e52ea2fffb9f4eaf86335eb7efd8a14af1",
      x"85e648d56d4e5079cbaeb8bfbd6d88567f2b74abe32b12a080920664029bd122",
      x"8caeb3d39d88dcc3b70c5b0a80131e27cc124dbe0a9bca001ce23ffea55a2a9f",
      x"1902e3d6a2f0c108745929012c89640464be6c762c14244c7d2c161797e73c2d",
      x"e75c9fa59d2b14dc560e8710dc7908cb2214599d6eee05bfa354dffb8189e4f2",
      x"c751aa72f1b2dcd8c157a857c5ecbf05e53caa234795ef5a6252d341cfb42fc0",
      x"a8b1459d2d0a700824ec5851b631570e78a690919caff74154e4908ee917c8a7",
      x"d105e3d38dfb7e052840fe008c90a782ffe7763de57f30413af7a315c932da33",
      x"6599576558bed85779efb3c2056afcdf16d2f86756f08ae339a11a919cc1cfee",
      x"164d374b32235fb2ad41f5c80065f122a308132340eb52d2bc5f2c1d10eea746",
      x"131225766587aba4365ccf586fd87e32eb0309caddb8b269917c508f219bb67e",
      x"a31334c18430fd56a41f0b2762571ae57ff41e84fff14a34c093bff84519f451",
      x"a3bdd286d13b77653b29a32bbd5c62ed27b9d2d27106fcbdec3e47927367c405",
      x"a6574b64d72014ab739db76424c7ed7137c00a2e86e3a7a4d5a79d33a3255f3e",
      x"82a05fbb94254c4f1f498281a9101ddedc21709c6bcd324eea415c718ae6ddfc",
      x"022372fc25e2cbd0afcff4110551a9f90de70e814d0ec910263e488766aaa7b2",
      x"cefcdd9554fb9c60ff98a802e1ec4e625e8b3508b036fca826b47fba6f488890",
      x"b09b3b71dee13124ee8f500f5b617788f5a7ffcb5d79483cff503641422d3a1d",
      x"ee3ba3974d0a285952a76d9de953fbf9ddf4ec9b520bd7f5a8a4a34fa88e8718",
      x"629bd8c815786f11eb07f1ee1a0b34ca23b75fa0af3d2d7ee2382e90ac17a3b1",
      x"e4d16141aca102bd161bf9621141d6e9cd6e011d0e9ba6846d2f453560e84cad",
      x"41655699ed6473ee3ad92c9c0157b3a558d2ce9fc15dc988475e319d18055ae5",
      x"65901c8d0401c53df915558136f10bf03f9bfd558ca17b1c3ec560cbcc1c0731",
      x"a52c94e8435a615eb911921cbeb6bb5cc0d8eb09782f504d326801626a5610e1",
      x"67a29a935f3621bc7dc15cde554f628e67bcf62a9ffb97b057b22caf6d1c428b",
      x"a544ec8509182dd38d625cf2b89b6abaa53c0d8fdd60687447ff8714933cf12f",
      x"f03c54c9cbdfc70f0803103c0456c0ee37b518c7be3fc8a1d82e5de313a6aed7",
      x"f541a546e9944c379ab2bb18414cf2c69d09329c00e096b7bcb3dcdfd34ccfab",
      x"5d045e02713a49a56a8fa322b77618278440418823343bf31f1a05543fcf0996",
      x"17f44d3f58ea331abf134113a6d1c8215e0a2308b96a56bc4b4fb4a8459bc0f5",
      x"16f7b9c37fc09239efdec81503321d7ff1b8d2981b0e1cbc251eb071439cfb4b",
      x"cc59a6042235b03a90be7b214ab714c1692de6ff6b536fd7927a74507fed15c9",
      x"ee9c5cc3002db1087c352457d8ad063bfa08c6c9ddc8283eff46a7f6f175aabf",
      x"34a7a4294a98ca5e0bb9f5311a3dcb079634776fa06e9242c486cd20958f57c7",
      x"27956fece4f8a7893cdfd18aa0646741f4e8796ba844fe80c7136255f7d0ce4b",
      x"d18c3eb101be72f49e55670913c144e0c5bfedf012d7feace40ef0b7b709867f",
      x"ebd99e5563cd05d2140f4593535802f6ae43e733b7d3704326ed301a3a675edc",
      x"fbb1c4a25070d484f7fd24de149933b2fa3682051123e7b357b30e3533903cd7",
      x"9505200da5924322a7a1b0fb9fa39e2b3db6ee9d449167fce661650cf9df611d",
      x"d219adc2e0680587b29c85dd189def5ab40fee381c74dbcc61fb7587f1328368",
      x"54a9afee492fbf5a0b1ce18edb75a4be346b30daafb5b926e62bd9d695a9fba8",
      x"0334106ac7aec6c0d4d7e404fe25a7920c96569b6bd0855aaec927588485a189",
      x"3673507f67eb407c895ac04af410b53265f9b4978b17f4adde8fcea164ae501e",
      x"73a5537157f97d67f65843299d2d0ac385d9be854923db751b37ded9d4947dc9",
      x"a81f07ceea2938c652243292201281f229c2ae59afbe22739134e15d5f81e04d",
      x"b79cb184059e0ea7c305fde47774efe19261eddd610e7546c446c71a62fa2fc2",
      x"82c545eb24ca78dbf66ecf1841a2d9708321bf8a66c0cb9e09642c9f738cf105",
      x"373c29f576b67ceb6246aa6f326a06509801bda5e65c4cccfdf09afa57a5826b",
      x"d5ce0e82889904c5affa5ba9983d78120e090cf01282a990ddfb43752c7a4118",
      x"36160cdb8bc52997b24851c06fd96e3a7cd2ac6014a8d5973b3dd7bf6b73a659",
      x"43286bac499c22a5208e27213cd08a3a47ab4f8dd8c236f59889cc7eeb8a441f",
      x"2dfe2c8479e83bdfb124e4a164041c13c983244a4cd23ac0b305f7736d2b20ab",
      x"822851a238f5c22e56ec0fe96ddd8cb08116116dadb51f5b83215a89d63bd4cf",
      x"09bf60c6d1e9925e540774c379a8bbfc16e34340a86d4ab98f3ecd1cf54ae2e4",
      x"ba925f6cecf87a3bac8479e4c8d276fc96e8d23a77cdae7b9ed23b751b580401",
      x"e6f2ff3770668dd5c4c13334d6bb1ef09bb4c9cfc392d366b9623eb37a91a7d3",
      x"2fe3c57bd561fa8a4fdc6cd24e66442e8b34bc1e2f495e7c57da56c373176be6",
      x"b03a3a5ca1fc356e5c7aad6dc14bae0378fb676510a875f36a7f1392a7240cd0",
      x"f73c7d09eec9c6f856ca184b69b669bc84eda93f728a597a02820d2ecb52a0ad",
      x"04654b38da87e428526d31ba1f2540cfb59bc3b348e0c726099098fefed1aee0",
      x"ba227b739cce02fca070d4b5a0189036e32d31d7f9087b33a12a8196cc3b84a8",
      x"a6072d69c5362c42135a7758352da171776de2934740443bc18231e1a66932ff",
      x"0af0520013921bf64d4756ee3a3f6c2b651d8bc46e0b131b1a02341dd1083b19",
      x"3067b7304dd1c18098cdbff427cadc15525d24052391c2b3b98584e6d1caad99",
      x"8bacf3a3e6f97036b593f6bc3ecc107f0830161c9629645673adff51e052d18c",
      x"d7a1a0c9dc61886659691122785860f3f01f42d42df3470c45207453a8c42232",
      x"6c797fff7d102dd00897dedc5ee7a142156915f8bb58f39549fe0e65fbb253fa",
      x"1c9d8758c88dec0835b5ce4aa6354a74f1802ff005b0a3f66a1bed4724406faa",
      x"7fbf61a979bdc21dc0ca7d6141a5a05fd8a020deda3f6536796832f43c6a3f49",
      x"77c81dca3cc7baeb286d7672109abb412efae546a3de1ccb9972f55728c96608",
      x"638b76da8ef427ffd3f163ca6d14da68cda7a4ae40d53c47676e371bb4f94ecf",
      x"ea54533efdfdb720d7398ecb9c6f9fde36f14e37d9229dfc994b32924f21f87b",
      x"ee319be3317608441ac62700e4be2c7d5edfb36308a8200006ac5032f0cd86a8",
      x"644b42dcf13d29013d9d2ef934aaadf0fec052c1f55f354d3a631f40f806421c",
      x"2cbb550cd992bbd150cf7c5e32b3af842c28113762625380e8447dc75fdaf9c3",
      x"9ae87965a55967f40a2f50225c51bc731055a649bc876caf9e9c4a127c39e394",
      x"5c38580fe5ea660f68ab72b1ad3abd5a3dbd4c42907d3c0370119153eb75c0c7",
      x"a0c096cc143e90c2cac431bba4716e10a2e974b20f60e7c8004f04b92d7acafc",
      x"a56e0bf27bd1a4dd08424f0801a8fd6c89604aaab2628d5e5bfecc309ce4a354",
      x"aa89bc76e83144a4dc10e88b5f28314807b8b6af0d266293927edac80b47f151",
      x"4101e24cadb30eebf4ddfd15a48be9357f2e010b1513def7f16c2502adf81869",
      x"13f9d480c7aa14ee95db237195e0098cccdc00bd2160facf6ac12b2278d61233",
      x"7fa6ced92280be042da4e3450fb9528052156497cf5e58ac47a391130df5ad0d",
      x"61e11ed24e95ccc993c00967ab9017df7b11375c24c029fa297cce1b32b40b99",
      x"2304cc3df11faaacce20330e9fc731a2098ad5047008402d4db5405068e3297e",
      x"6c5c371800b0f5a3170ebaef734aa0d9cdf60a25734ac1ca649991045cbb1802",
      x"a8c322f5aa696a1b2c57009244fdbf30260104337d8580cb33431c34544a94f0",
      x"e325deab8e32f167371665e7f525f8d17f0b94005009f52dec3c0a2069c3b63f",
      x"d076c6e020e3871dbd0cf182936a2ce53ae7f7570de78685c3c417a6a2f88c03",
      x"84abf3c2edfb04f7ea8a1076180812eb0e408b5d47f2565cd564eb4912570b20",
      x"83366b970698a1939edf238b7c399966b354a91c787be454ebd4eabe3de83811",
      x"cd030e8724fd29a301b99ef4ddf78469a7490a54e76349646004cd46a8288869",
      x"09525876e829485ebce3f487d76ef71a3a527606bc5485b80b8725705fb551f0",
      x"a537c7c29d6c25dc8b6bd3f1809ea19c6f0591f2cf6b1411007d5d863f08d532",
      x"f7e7f9433d67a96e0b5ef84b7c8f0c09b271ede5574736524f2eb85caa5bbe56",
      x"7333941aa592ada42f8988e15be807ccb78df2e07df7e4ca151620887503ff80",
      x"e81815093dd1bb10109a101e99d024314dd861f4f9f3489901664c048edbf99c",
      x"28c4becadbc00ba518f138fb386b20b3c080aa132e8fb4a8df265a7f8dc095e3",
      x"88a929a53db738c8e991cdce635313a13ebcc3902354b7fc3988531062ada78a",
      x"6cd0821dd8239bce83dc2d4d734addae8772687beb4870c5a73d335e43b6349e",
      x"c8b3652581033ffef17a4946c010b7df2617864edbc936671f686daaea0ea4df",
      x"5b3ad4960cf5882a02a09e3295d7197990f24cada5d058ba8af46b1d186a0bf4",
      x"da726adcd46460512127ae682813514b4f02a342b85316dedc4c8670d482bc72",
      x"4cda695430149574fe42187216e20a123aec599fabf7cafa3685dc5dba049f80",
      x"c2f03a0b406ed7d04b809eae612e6641e48e5c9336b7aa8636e545ba1ee0341c",
      x"6df82958b900210a113273d6bb8cc3e2be1e5b7a1ea42a4d86c9754b399107c6",
      x"c1e058136c3133fad3945f0688fe5a2d6922886165d0eb23af93f8d5f7237c89",
      x"78d317b5dadca739d88954b122610deba6bbb238f25f7c97595a025f7a584906",
      x"22f452f2ac1618529ab9564d23fc75ed8843152fd6e61ac6c1c0086d03c7a9ef",
      x"845215a8bffd71dc07a65d4c31d3e9881b9c353d1433543965a81f6098cb5ba7",
      x"7641f5149e9c34c7efb9845a81a366a0000c0b188ec7c4c29905f8b8e5491604",
      x"cfc7ab3272faeaa333ec14391e7390c913eb91f12283070162d0fbe429a722c5",
      x"8d0ce57326450342993f7fcc1d2e8a3eb41c0a1a5984682031df7bd7910577d5",
      x"6e79105fe99ca4b20467284d2e1dbc142659b31d248530e479d567a8bfe354fb",
      x"f07bfeb17f47ff8778ee225079cc07d2df5aa463765d1020e11f24619f5f1873",
      x"69c4ce4dc5d2c6cdb5a40c2c485eefa7f7b18f66bcc03a5e813753431c2f2398",
      x"af8d8ff3c80f7acb0ebc2f00ee8191b2e314eac70e3371601e17c4b56774d796",
      x"51d3f6bfaf6880025319b14abf16a30dba78d30bebb5f140d76886a9ab5c426b",
      x"dfb01888022707ab4ac07dfbc4423d939ca7feff266444f6e6585d9b08ce2c18",
      x"92fcf2e5a98961c5b9a6776d5fcd36e3c65b7577f19cedbfd4b6e6b9ea48d529",
      x"1eab9fd19b52f2a6847a120f35042d3f7879af29c5915d4962c3e3dd56726784",
      x"d7edbd9c9aa6fa1af5e71f991e56cd3c208412572fe2504e769bbcb49ce3c22b",
      x"398c2f5d3d6506acb8177675980c7f386ffa87f8cc2c94e17118d68d38ec844f",
      x"c709e341ae8650c09647fb8d8f999b77af0d3b2fd0efc3dfcc6684b68777067e",
      x"5278c7a742a48ecf91e10706a89ae44fd9e54fc2618716dd4d7b8387f3be7172",
      x"3e27353af26f20f1078b6f48b152819d034e96413ab88ea491bb78ca9099b2a6",
      x"53696fe05c59eccc81b79d222260629577e09897ac010e6a7ac2de134d190eb4",
      x"817f62d678eb2ba4c57b3e28bdd2d965d5dee07a2bf7ae799a6e3f2d64c3de39",
      x"2efe26588b54b536eda538fa78af178f98574a394040d6006d706ca15698479f",
      x"ad6c7040482b34567ddefca4a37bb0a5f8cf4ed72e331556eff514d8bcb13dc8",
      x"58b3d5014a44b167224d82b8d1abbd574b6b4829dc9733a93fe4ba72977d513d",
      x"5e305f86f738be07016af27a7e5f5baa28c85edff966a640b2183535ab353c96",
      x"127737c38be55aa4c39caadedd751e223c82c19eee6c5164554be4f509674658",
      x"d9822cc9b6ef7f821af5121c93a7dc85860a140f504ca01f4633b1b2ac15b5af",
      x"4ce716d4328e19a2d89ab08e9246ac174283a51d817e1865548e73eb38df4a52",
      x"650dbb4d6d691697efcece28efaff6a1116777ffefd8a61cc9834eef2f09d5fb",
      x"95bf76a0f43b308246ab05c4ef4f8f2e71b33f08b89d83ab0a7138cc25f22459",
      x"55a1cebff524499db643f874d759ea8fddfa8c38df4dfb00d9622392d1c49d2c",
      x"65fe27129f05615d9defa7297fd7452ac1b7a949266c329dc51ddb815bcf5b32",
      x"7c93fc514fa80a0670df3d97bf0c2e72bb0dc602cbdf76f5d6006a49a155b418",
      x"d8edf7d36d59ab7299a8b8ecb5eff63b951265268b85a16f3424abb58a62ba06",
      x"952b4d6258738fafd72831fbd042b7f7b6fba45f49ff96c398255b5de8a20b0a",
      x"97a2898712e53629e31a20206cc82c8fbd01ad00804db30c3b589f0c28feb50a",
      x"900772b3eda0496158b0c7ec6d73e4c323ad7f047586b7f019b9ae8def229f66",
      x"81e976119607a69772094b1786e487db729a7f67af6e426cfe12c57d9c972c0f",
      x"8c084aff910e8c9ed214837c3d5abd21f8d4b7a4c24179257bd44b82853e0504",
      x"749427a43d20afd45faa3b3a0fad5e64d2ba3ced38f0c229944ab1fb92a94db4",
      x"c550563a033d6e3f474fd5ceff1d1f4cf3541abcc53783720ca45799b3d32b31",
      x"a79fe56587c7dc5682ef3cac904838db5fa724ad26bd33a9b41341b8d7b2a344",
      x"675627e247074234a9edead0b201d4bd74a19b62efec2475f62e8117a1e40cdc",
      x"260f0cea1049c3899833c641f5921818b967830aeda4748f812c23db53c25925",
      x"fa7ad05020184c980d0f72f642887ec26d7f1bd638cbd8b15193b4ce0225dbf6",
      x"2f10814f01426bc06bc0b00d706865056d2b33f99ea983eaf9ec7b263d8341f6",
      x"61e1ccbaa139019878fa3a11573585847b0239728e923c7b19ac6d715acf8757",
      x"d5f87747e7d995fc4bd03f7fb9b58a2044bad46f8dc623588a7d82e29a20ad68",
      x"56dd30edc16c4ecd607c985e8ae228a37c2eb298229b42b2edc31e7a0a0e9a97",
      x"ab95e38197e4d9062d889e01d7e236025616b147a97382cc57b2386eb468da01",
      x"da913457cc0db2778d282f2e0d7ae2fad551f85515f0fe0176d59024996c17ef",
      x"d4391f53425a86c9c04d9e177874323aa3f237fcd2e01d13b3ceb7adc94bc757",
      x"f683a2afabdbb6aa4567676360fa3f5f192340fb4027a821d52c072f1a9e0717",
      x"66d3a002d9026ebac8261a9683998744f96214ae43cfec07992db410af6d4c98",
      x"73b741d165efd0c8d435072027a49b4a6cfc35deed927487553bf339a842428d",
      x"65b6fde18decafce57a6186de251f663cbaafc6c6e6bb7bfe8abea4e43b7dcc2",
      x"bf6f20bea2f61b606d23869c42d4df37ff8fb5dcdc15103b82be023e05f121cf",
      x"0b2ad2d9b6cb2fa73dda692ea0d1b673513c8bb65ccb58a02679adc71bc883a1",
      x"880e892d3c61772f66ef995c7a71509155851b29dd84bdcd17c2d02e5da6be5d",
      x"0703c3c08d0067e98113e469b0a9c887ab45533d6a98bb317003ea85df8f8c73",
      x"b5daddbe1a45912865c88d6ff7938e4c564e5b6aa46d9f1ea822c90126760861",
      x"e1fe0e96828d3ec81bc80ee4472b9a8c9e05bfe563be435349334c2b8e18f05f",
      x"a24f09468333dfd66b87d707d8ff57513a218cccddb789d6ffb16bd9815c0c98",
      x"31f7641e04f574a7745129bc8ab06739d97d839d7a2bcfbe52f5a5c1d9c376cd",
      x"d39d658bd47da9576d51a105e37c7d283b96877298e95327373c46ae904fded7",
      x"c35ec1de4f50cefb480f437fecb9396de920c25ed3b904cfb52a4d731b426231",
      x"8595e21d6d8b3b71acd62cf7104db0fba86c0856f580d5fe3deb30ecfe0091e1",
      x"aacb53401c8838e6b6d48c3f672f1535534236052edde5e7512409c5d9e371b7",
      x"9216e90ddaf446df3287e325c3088637a55798931cdf88ae2b4d215ce1dc58d2",
      x"dbf4fb918035d3686f232bbc2239aafe591b512e6a71470f31a83674d66b5fcc",
      x"6557f31684cd6aa9a858573aaec3b1e80adf02c2b72d5c0e3bad561b447566cd",
      x"d4d251d7550162ca60dc67b480f59693804e181928b9099cfedc490c84d55572",
      x"47a107f02b074cca3e0473bb45f93715ac01ef80559cdfe0e713d8c44acb6862",
      x"230d45e7541cfaf160110a162b16b5e821a0af5f9f50117341cfa43900299bf0",
      x"db5c096f71ef2340bdd9473733516858f0f078f37527a16e4e32f1ebf8c6226f",
      x"59f7caf25ce714d76dfd9c5a172f5f68a1c0fad95516a1141b803e3cde8091eb",
      x"6a0d2d42b79b9108fbb935d0044bd7e4704fd12285eb32fb98ff4af23ed54788",
      x"6944727f41c746ddc3f16bfdffee6e4edefc1c7ac9dddce3f84aeda1c314439e",
      x"6c7d3141bd96e2271d8f31edbfab44791b8d7ffebfca087f2fc3a8339cc5424d",
      x"6d65483cd2b1d55a035a36e740da0d7fcf1df9fc18f70c2055e82fc3daed27cc",
      x"c88fc65c7539266b318d55b0c4e7fbf148a4cbe3be250bc7ae675fd4f057c1ef",
      x"284e16d2211a1d5109d52c102721f30bee827ff89ee19bfdf8898b6f03e837f5",
      x"ddd3043262f4d6bdc85ac41fc818a7fc2d2cb703d5dc34d0c066f0b513a7d503",
      x"4e05d89493dfd0d3f9bc75a954c0823ff7565811a3b2052002fe132c8befeefb",
      x"a52a83117b70e81c419dd44dcfdab029020bfb10b05f968f2dc0b22419163a96",
      x"ab9731be37e5ba0498ed2fa3203e2c5dd88b77b663e75563c534c60711569680",
      x"0735efe52924f592aac323e59312ae6d95855fef31893730d6175024f05d91ad",
      x"f1e6faa7c50bbf5ed116222a8161cc05cb2318e962f9f11ce72d113c7d359633",
      x"af584c093d9a2f96635ea6ed9c63454931dd1d7cb7d38db58b350d9a5a1800fd",
      x"453dce3398e136ecd3072e413e30fc8e2488766428b78dc64cca277543289f1e",
      x"d57b9047236f122972395a5b5c12a837b34d84e31fa9604c4308626e149ec0ac",
      x"68bf44c7d188d40344efcea3130acd94bf9b8c467d162a3717f940af30969860",
      x"b9f5c367f1ad58ca81cdadd90d3e36f106ea1d20c2e43cce3bc2fd828e6ef397",
      x"349acf0419237a71895bfe39f2e20a8598b83a1d953031e5ee630f5c0ec65f86",
      x"178d13e90fd8c813a892503010bd15ede13a5b067fd80453f7e312d93f81f4a1",
      x"95d8d6591b2840e726f97d3d67e35b1204bb847095040878ecc813a8eda7054e",
      x"cb8e50f7dd83c783e18d87fc8734cb4bf18c2268d358ce05b26d93174775a24b",
      x"796c0f6b7d449c3f4008191869467b6bfa17acd9a0573cbc290e807eeac3d2c9",
      x"4b115b8fe21a5bf4c4ae615127748b21558159761b99d6f3b21d72950e14cdf3",
      x"582489aa4cb2b0c755d7dbe89ba90a920c9f094a79ad9df770a2bd2db62c148e",
      x"ae84e0bda612080796716cec305deef8f6c8d428135b95126ae5620083206a9f",
      x"d5411b072f5a84bef92c2b7147069932fa83e8048ff352f620d0040b47f323de",
      x"48197df08077232b6852c241c9d947545b585d173c23b6f26b1e9bdca99c0595",
      x"0a77b95cc6fee3d261eb012878e7cdf98892a7ff096b642e9c33e3aa9b5763bc",
      x"70eefd4c938a202e0958cb5bc771a09a5c5dc36b118e5e71c9549d2da1771e1f",
      x"bad0ea55994dc76e847d245270225d842fb99a857d1636ae8e8c94681bbe8118",
      x"8098aa197b221ce69c1fbb66a066317007552eb43c24e6d5d48863fbab79d206",
      x"45ff4f40a59005a6c3dd27ae4cebea300b85f17cfd84e9140f36d08a637ea63d",
      x"822a8ab85f0ac3b957ec32e6890ff922bfe59db7e3d06ef8a8371a6d33f9c8e3",
      x"457c11bc0457936055519cbf954bec593f1b93a0425b90fb7da00f0f52e69352",
      x"2dc4f6b85e756fa04ff0f8c5845133227c795e3f473b96870c3793f7ca70fc98",
      x"a38181084fb8365ceef237d6e41d8582ebe60e1bc1c7bcd0e09155610f2993b1",
      x"0ecdee65640e567c611aaeff6e12ad1fe48f7e94e9004a77975df52f4473d0a3",
      x"b139ef543d9d55bc44a8897ccaff87c2467803e05f4dbe1c3122ee0f74c05451",
      x"c10b8952581f8ebfcb250c69edab7b859e83f171c534f0713738339c3773fa9a",
      x"e29f6deaaa4568056748f8ed7cead518d038bb46367a51357a987ad4e6774e9c",
      x"7976ed00571c7119ea9569d3d836993a3b8ef2b70175bfd3992bd8b182c751dd",
      x"a307220b7c7ec7e7bcadc15c48e729b19915443fdbaf0e84e9789bd7d1ab8c49",
      x"6b130bd75ed335d697c48b1f810ce4ec2409e77944f9371452bceaa2835fed87",
      x"7969bbd93b9e2c60030b0ed59654b39d18f45cdd470cca861d0e7af88e4a85cd",
      x"2c1f7e193f5441a640d3b12b5afa9f52967dcbd417b5cf2e7bebd329c66e8c9d",
      x"2a81cf99825117fbb3fd902ad8893ca4ce6b8432012ff082fdca2a9dedfb8215",
      x"3567168c4fd53d33e685fd20a0d881b917cbb5a67a0be8a9430c82d96dfc127c",
      x"e8c8fd3f502d57a9dbbacff46339d2140dca3a413180d5d8429b8c50728d1a00",
      x"ddeebb756a29e88f5de38ccac1266c6a00e9dacacbac5246dabed765d214fe1a",
      x"70d0c4918e6ffe8ce557bad515cb0f24e0b8088d9f07d55d6700ec1ad6ef29f8",
      x"c46c9db1e2e3e8befe110747d5f7ce1bee3bc5151efa3ca5da8b9ce5ed462447",
      x"e18b4953f7fac7089462c95fe4b86551690f93effb9fc8717a9953ee802bfbb9",
      x"5f3c7618d04b457224ed4395a8f715c8752c43e82ffe0a392fb79e208dd14429",
      x"3b261bf3a95dae6f837ea300760f437e036cec36de45286c2387c68e1c874be5",
      x"f8dadab6224d6ae33cbdb7a1fe5a2fe50803238a1addd61e979240b3e021584d",
      x"0c2eb66e5fef963d471ec2c666dae753b48dba2b78f0ee74451ac1125ee68102",
      x"8f13a7ccc2ce5be802fafbecde01f7271a41cc3a5ab658a8d305e670780f928c",
      x"9ad0196bf14ee958f3736ea1384cbdeb127ee83012da696f822532d7931e77e9",
      x"8c1bbd49b56a8d7b30bcf38101543ce9a470daafc4f986ce3c649e7b62789eed",
      x"e0f5a8f269fa477a0d1f9a64f4da499c937a5b1becd082f5a9db4053a5f0377b",
      x"8ec02b6a32555141b568302ec8a57fdd98ab1a312922f565bf7cd6d31f029605",
      x"a7451e178b01eb17146e462bf0e3a0d4f0f2067ab3f0c1bded7a1d7737c90983",
      x"6e32c29bc593c3ad0b5c3b26f67733899ed3e1f0f76484647e7d9899dec8816b",
      x"89628edb38f3bc2a449d33fd28f9311d03daf76236abadaaed6f9103a79b29a9"
    ),
    (
      x"46ce4e86485054e862227433db193a33fc5e36928959e12eaafa977edd97ab5c",
      x"e288cd2204cdddb02984e999e2d6cf3ac94a4978e69748c833ca0e5dce39e6ae",
      x"930b1b83684f0b20539e02c506e0aea16daed58c0ce0a176a144f6cadf7e5f0d",
      x"fbe4c64075a468d7337a50e84f08c3cc81db480483d7e5f14150b1e2a06ebb7f",
      x"69442ea3faa5e15780233a4a54d37a8f0df2c82ec1139f329e8742383bfb4744",
      x"2f5caa211e44f2f9779711f0d7f320d8469d1701e94f73f501670d3e930d75e2",
      x"1b1f76a23161415c43dfe837302d74b241c0818be9230a0a5e0e2a5ae2c34559",
      x"9f0bf1f337d5232d24a3b690fa9c450f2c2deb56055d13c4b875296ef1c047e9",
      x"fb3366e560c3ea98804e856a2ef3f596fb88ce57e8d922bfe16f8ea63c6a1bc7",
      x"91eb8d07ea8bfba2597ee195a5dfd891f2b7b9d3c8f43178e6e14ba379d9e86f",
      x"5f757cd7d76bb92a89798ed56f8cff349e348a729c124371da5d67be48bd6ec0",
      x"a3046bfd82ac638b6e051310d23ba4a73a58d77ba918512ead1c18b5eef28df3",
      x"dd610812a9303f307fc9e72150983f2f77686f33e63095e881ae1ee18c1b98df",
      x"f49291c008d2199cc19edec20d88dfa5e498036b4841cc76233bd27ca5241fd1",
      x"e8168454c302652d3d3acbe35e0456d0952a9bafba7de14b93fe600f7208560a",
      x"401506178c55e670eb783e32fd579d0649d0d34d1df2c83f9319d033cd6ae79b",
      x"193809010a9b390f556c969d9f43c0377a3532f3f1af1a7cfe2faef567584e84",
      x"292c610657d75c78e569d2708b4ed907edf533897c96c6e3c4309303623be98b",
      x"2c81f4c8f8a98da5e1d8a117fa17601605a960df9f63bc06cff5d09eebd974b1",
      x"81d7db8dda7834ac6cb1f24f1f94c2888cf440e0ed8f99f8394cef42e34eae1a",
      x"55b0a0e5c3ae1fe1014cf4fa32acb4562ec1546f0d1e48ca6d76ae709d567547",
      x"d1fe5a8a15fab98fcc1b70aaea119d7f19eb45ae6248852df0575fe24a0b397f",
      x"645b12c3bfb140e3d54d821856218d0ccbc84822d9e4edccba08c7cf5367fd3c",
      x"aff88f6f4a35289ff2f8005113d2ceb3d1b7370d6728513524a5d1d62d597499",
      x"d348972d3ee1a0df4ddf62122562a170935dd5903e31b76e2b6d42bc23f6ca7d",
      x"c4d4a35107af4601bb641581510a6e7014f2f76b696fd5d393a0c0fe38481057",
      x"187714e616af69499e1c42de1354f3b2eabcf366adb5b46409a0af6aa3903bd9",
      x"1f6768655ea6a5be67bdddf1629bc489050554089e3ee06404a47afab79a96a9",
      x"a7c96a6bbbbc2a26c4d53789cbf2cf832a9cbb6b732d089c712c91492c798032",
      x"74638cb9c29ee5f8dd79a795326862ec3e7387bf660f2a4c83b7b5be503cffbb",
      x"ec0949c1a8a2ee8708b006d646ec56938adbef0bbede0cdf38b567a33d3f0d25",
      x"b19d2e89605bf89e45c1091667041c3f0bee2b384567da411b0772c6b68167c5",
      x"824c76218828a98b402c1a1973295eb92a1e6a707d63848c5a7701b280616388",
      x"4aaf9e5ee57879e75a00e6f86aa8916942a3e4125216542159aa263e7e5c3d91",
      x"451b4113bc88c983ee85232d0cc36cb025f2bd30b987a1813269d9b0c7d27776",
      x"3f1b2b110957407567f7918f737e5f846ad7f1bf81bbc10219ed82b3281107e8",
      x"1f45547068ce0ebda36ef4575cbc6a41a561aad72e2d0eab9e87087c8064bb4e",
      x"ca838c75ea64740b19f5b202c3f42cf28789b3f3ae784b4b9ec1a944f7251c26",
      x"00015e8cc26f7eeb3bab163a5f3d7d4b128aedaee718448727ae22967f87c05b",
      x"c4f572791da3c9d198dc274672808b9ff9e6e98d968350253fa5c09fc7d18b41",
      x"84bc4b578bd87f267ad59ed4f067bc619d83a78758c82dd993c75ed5bb4f222f",
      x"9bf7847a723e6b4fbc0924bb8ade4af8d4743bbf805d3792994ba8a2a21620b7",
      x"23a80ee1e95cfccf0bd16e8cfa3ca67759c06fd28b46ce1fd97554a56c07b448",
      x"8747d6e0b7e7bd55976cd04822655e033081adff60b6e0157029b4e26ad6fca1",
      x"7f121a0eb5e38f83444fef8bc35825130a9d9f3d1e4257c61dededed694cbca5",
      x"74bd1a6faf8ded88a1c03d34f7b9e6376f759b915585408e1b51696d83ba19c3",
      x"ab358c0908c0aefe074842e16b5a0a9d9c54d6d4b920c26191786be0e44f213a",
      x"35618a37f438b6f0aa0c682a53aed679c098d823056511328c103e8dc9d352e2",
      x"d3c1edf6ffb85c60813de15053855b20b46b8263c1a1df74f547e0a0ebd683bd",
      x"629f01fdd0e245357b23199f3f66d321e93e5201d63edae1ff9acc8c96542dc4",
      x"e91a61c17c65239ba80e4a511e2608cc8ab2158139a1a3fbe8c37efe9da03ca6",
      x"99e608932c8fedac878c2c0b66ff8a6686e661f92e20b14321816d24f5dcada5",
      x"195c266695a205412be00861c17bdb66bdecb3fb3e2f3384e16e5a368091a4f2",
      x"a7204005d7c30347e702df47fa3c24a6235baad7d3089021d359c5e9f71b821a",
      x"98182f985a13b530018b323a079e29df6b1203d88ad74de9c5aa7ddbb03e5376",
      x"a5f5aaddd86f3dae605afaa9389f541e08971e62400321f8961e884d4755f98d",
      x"30bcafe93b0e7928f225689af3c3bc905c0e6640aec77a942cba757a63244d68",
      x"42aa03f3f37db29718959fb2c818b30cf2944f1ee9016a1f12979af735f87fb9",
      x"c3e3acd3371ec88e34f6a7be1ec325343e635ddc7725a61c2bd541fe08a34458",
      x"adac05e7a5e4aaf634f5d2e06024dc204bd384be9d8ec55d60af9ecddea3db53",
      x"7f2353e239452d81d2288fc055a7d1c3a83cbd78ad6aab6b2cbae1ae3bc0dd2e",
      x"449a7360e98837b510ba4b72aace8aeba8e60a5d8eed17566951f6b657ad36fd",
      x"38a2c02a18df52d5a37c00430ba2649166f30440f103dc4e2131e6f933110757",
      x"d6a8599b2046fbb81f5919b61d9076420ba3d43ab387101b7ce6ab232badff9c",
      x"7adde850b176d24297336a194695ab9a0bbf3230b3f989e41bd4d90aa04beb6a",
      x"decef3ed981b64661ae3bb2413cdb0d084ee129f6367324081452774aa4c1b0a",
      x"9b52e43530c17b369af80b5f58966d7877da1d4ba08379f4905a6cbe8f00590b",
      x"101967c39e2dbeef591202ed6578fddaa1c17b897586bd124593e680f912861f",
      x"64425a0acc4ca82d6c135e43a4de503c1a55fb905a30f0de0cbbe59ed37daa91",
      x"3bdc9fb120a04c155266a6b6c7b59c4a38cd9b0b76ba6447f999d31acc5d535e",
      x"08c2703398dd461c68fc68572ed99a5120b2d810b0a2b1dbc7de6c94f7b31f7c",
      x"0c79b758f4f0896cae4270553e5682e0fb2f6cdb4564013e3a8652df6d148353",
      x"139bce61624d5d085b2e4692ac44256beb310c74d7348070dd41cde3c5169118",
      x"d71c9c89190444dc4d851ac14db0059a0e5ef1402eeeb025c8d48dde5e9566ac",
      x"7506591063bfa93e7606309e84a0e353cbaf33afb50407e0ac372ae00c771b95",
      x"9b160ea72ec727868899257c3606d0f15c33561aa274bbc4efb21f22ef1e4b1c",
      x"53336ed5bb30acd5c5cbd58ccfb4093d420026fe7921fd9887e26cb178504f4e",
      x"91329a346da381c57038d297467ecf9cf1c6b430699ae42b2276a7cd5bb32d5c",
      x"eb7c18fcb6721105cb97c9ca7f001dce78c2321285e7bbf260d675890ae1bbb5",
      x"d4e44e561693b9398e13fdcc38a825972c28eb5ac71c740f2f3c5c4343ec0dc3",
      x"ef32d0f9544043c25d2a619a3af0638dbf8e413aa79e59ae135bfca38bc0b8b6",
      x"f9b6b15fbb6148049e63d32fefbd0a26553381913f89343bcd6a48cddf707423",
      x"60481c8ef810b0b116f78575ae34c3522e8ec70764820c5ce9d1869cbd51ed45",
      x"1aa144bc4c8299f0be4e30024f95619802ad2cc51c904da8a3611c6c7df0a37b",
      x"67c141253f1786686eee1bd394d395befa7aa8b9acc4351036a7373785f7a573",
      x"c56c54ae7038ea77c793a2477811717c83e464e949b744ae4c32d8070294fb79",
      x"f6e014e4f8b05f579bc733b33c1565b681abcce365c3ee78db69166984f1134b",
      x"6ceb018a0410019e01e42f7db5a49a4486ec53139d7cf744ca72c97bc04bd36d",
      x"9021778e01f8adcbfd189e09dba496841e971f40d3bba7c498f6b8e61d3f7211",
      x"8ca7a0a50f57ed636b209b6edea66037fdce81aededb833190896f79d30bb56f",
      x"e7e98039e64fc4b1f83898490dbb22aa4a96e375079c8f931300af43634e41dd",
      x"eaa3580ffade491955c28038a39d825172d3eca7542c0da656ec2657e51e507c",
      x"9e740e235f1afb1d386ec7c0b295299c039b9dda1b1b1f4dddf358b9c2394d73",
      x"9d21a9dc8f8657cf1711ca65a54fca9e1d806bda07e0885dd31e2619b8eb69fd",
      x"c0eb27fc529903d212ad82808d89a6b610b1a53de03cacae80d257f12e7f86ea",
      x"0a7e63faa82e8a58af6fa0e5787c286fbc9f7138f6e04d2aa523d9308331cfa4",
      x"1d5934b5d7920e6c8fbb6722438d1d969d0c6fc3e50329bc69ad8c3341b63871",
      x"e9cdc04f3ad9a3bdd8580fe6bc7725f883dcaba7d914953bdbe8f7b12c37c994",
      x"8c3b364a5a0e99c976d99a7c03f56d6dfc4c881174072682f220e53ccf68e906",
      x"ad20d92c9b088f668c18176baa2c9b381f57a28458b22205a4e0b50f7bc85e3c",
      x"c539816946c7190eebd86a551ef4b5841236fb9530448873ba869dd90bdc2a38",
      x"f9248691b57f6a9b34074118beeeec861f836a689af44d6b256ba5dfdfe2dbfc",
      x"4d76a57c51430803651e0f8f1890252b4fd9272fcf76a84dc1dd8257a6ec1fd5",
      x"11d6de302ba6665a5daa06b8527ccc8825c8da39ebd9b4d9e1a9cf2af40c2544",
      x"c2bddf86d317e641ebb4d03aca9541e7ab8366d30073154833e3a7785bca13bf",
      x"b1bcefc578dccab331205d110c23f64be45a00058a7ef3b3aacfd42c7c495dbf",
      x"7b72e68cea9d24c236079fe4639b0d88633332750e6fc45828f20f95aaf93844",
      x"b55afa1590101e5832d19004776e259d0e5edbcc51a34aa70026a6674980b845",
      x"d0e5fdc7c20b5ebd19d0232e3c882e284c29320433759a588d554b1cac31580a",
      x"c042a3ec33e09b03b08ba05f5da60ed19d189adde65a0bfe6284e4ed3c943520",
      x"78bb61f4cca4266149b43b3dcbb52ae0c82fab82d9da63f8a66ac6ff84ed3fa9",
      x"88eaddd586ad5de75088c97ef4ead0b4a565483382a2b996967cbdb3a0ce1993",
      x"baaae1f03b93e495b46498f6702f5396fc7f22b68dd7675d533409f4d393e92f",
      x"a80462d63041801b37db10bf224ed5ef0285a9cb1fad63991a494152f51fc7a1",
      x"308feb330dd49654dede639bf5e372f80c6608c6ad2a297aa08ec3cd7ae5f354",
      x"dcbbc805ae2d6ec2ac7975fbe3394eff61d561d773c022acbaeed049568b2292",
      x"59605b9ebbab9a4aab4850ac69d87986b6e659bcc4659d20bb55bd2103713a8d",
      x"46bdac5a34725b63e3ec29b1eb5b36d979e5343a8c99298d67be3b2a386b9d45",
      x"5e4c711ae2c0826c6b5badb21ce0f546f32289bee9df10841dede1c936edc4d0",
      x"dc1e2f1a0bdc981e1ed59a441e0fdb012631ab8dcf490dbc40e3b96cdc8bd66a",
      x"7a241951c49416b4ccbf43b4a790836ccb843303692cfe8a71f539954a01da67",
      x"ab61174101b33b050707569bd1eea96e14f2a41863cb98851f842cb6c28e6b08",
      x"2401aeb4c6e9f8ea6ea70e51dc9c37605a0fe6f7b33c0faece104c6d65f83e91",
      x"99924572844ac057e1be9155f3dd4f4770f21f0c132faba9edf3ec5898da6c67",
      x"dc873b548ceae03a6d3a53f6493e63bc979e70b4e2bb5b915c101f88ae7b3a6f",
      x"c0bf7bd5ca4ffd6d889de6b64b2fb611f128ca2e85a703a7154d839ccc6b8e42",
      x"da476afa8569b30f015e3ad62eb63b20bd3da8b94490c08dd49fbeeb86e5be36",
      x"d176d6148a85d16dc10c05d868df3a283fdff73de4dda20bf4df8e2f4f6f17c4",
      x"8f9e0004313c39a77d023e2ca04ec66c3a168c89d7bc837a514610efad4738fe",
      x"62183425d5e32821e61b020b7173ca7ced9a152f5fb19eb1451402fc8bba4c73",
      x"2dc10169b6ce86e8f3dda05304b8753f658afa2753678e6d7dd6afb11ea4ac7d",
      x"fe58e5a7a14eaa84418dd1cbaee583208dfdadc5cad983d9838905529b92acdd",
      x"7099dbb9451f228608f04285cf89043ae70af8bd5a4c7dc195bad79173462775",
      x"cac71b6a15965ea14ea024a893b4f8c09637a1b93d754db1b444eebb5ae7c770",
      x"797cfaa8c062674b592d0eeb5a87cad4e691e3ac7ffbf06611e06886e1faff4e",
      x"25d288f8c6de97386c2fae24dae10a8aa1988fea90b71c3f04efda45558949fe",
      x"608cf26a1852713b976c1ef305e7c0f8a0495df1b98be895ddca111e8d766661",
      x"100d073a480dabdfbde7cd8f137170c53a6170955dcf5db0f421f0021d87a5d4",
      x"4df4f89b03beb3a72bc21a171f40b1c4f22e881b38cfffa35588b48b337a5568",
      x"4b81c3ca30f0217747ec8bdb6512e1c1a35107ab99448621f1295b267b5d0bb6",
      x"63b198adb2b6f95994f5063218fd6753f4bb241403c13a58f8ec3d4fd0bcb0e4",
      x"aaa2a4725bd20ce337ab387242cca5bbec7db1243417afb8ecfbce07b16ae714",
      x"44fe4e6ff11b9d24c01daf4864eed50e1089b6cd125950122ed5ce94dc98d4d6",
      x"5d64f89547ec42e1b892f43b4295a09c5aba6e8050883c310568764d6b8112c0",
      x"479e34e128179871c6f6f673d0a808f65083174d1a3b4b0b6398cf2c08607973",
      x"00a5047befe9e94d825a1d157b4dcd83c601033186190fda9aba53df0df9afe0",
      x"a731fbb87caa42278f0573d41adfc8336f3f273bc0d11ac6a79d6c0dbb20302f",
      x"eb8857d2f450a7aa958b04bbcaba359de58538e68e6b68f4abc0364ab6f0f2bd",
      x"6f9abe68ff3753d595c6c4e70041efe4f21b9e6a2f2b27b78b352b4073d3393e",
      x"c4e5921d11cab6da3a7904a2d06f60b103bf7734f5dba4e306adebbe51f22e09",
      x"ee0070895607a08a1c339a6728ac1423df26942ba900d73a9856702151b1d222",
      x"41114c8a597b8a8e75a8cf10cffac64f08f753fdda71ada140783402bcd034ca",
      x"9a103e02331b0133d4f24d4656ddd27c76f3d5f556db2dc2a7c7563e5f227b7f",
      x"1754bfd2e3085fee987f523f79d299d4bf78ae1eb8a9071694d962ad7a8b8a92",
      x"74dc2cb04d3774ca5b4b00b134ecdbf7f7d90d0c4c2747508d1f674625cae8c7",
      x"06ccf90f159d406333abc788ff45d80d381cdcd0721253f13abf1fd43eb75ed7",
      x"29c995e88bf417a90228960f148487f2d93b4c2dcc4771897fc65561739a5d9b",
      x"5480e7b906d42b527430d22c383b044b0c9eeb34b38bbdd7c1e0932a515016f7",
      x"3729c79f46f6b8110567fb4e11bd64ae5cb3e036132f845c720a8b6f96df2a74",
      x"414f5afb69f8f35fa9ef1c24ee893e83f6e9d983544a46062210e51275f46458",
      x"4b0b1ee86a1c8e0c266b86e89c2abf44317a6c242aef66cb45d5ec15c51040a3",
      x"25822d7ff967eb1e76a23629a1689cafafca0458fe64e68e1845af6e4cc41c58",
      x"01c723dbf155fa622ee94dbc72c03118c71362e97e808a2d3809db0ec981638b",
      x"e71f27950a828f5ed595a92ecd66126ada7e5225597973d18315e0704dc34a3d",
      x"86cbf26c3c4eeed16480f4d3c2977fbd0e4aae50b3398c31792e2cd126bdec6e",
      x"72f0b69a877e342414a1cdccabbc65cea4ba64b345054c0adb33d8b8e1924dc1",
      x"73be58280846d04539dd2eec6ece05fbbb0d8c6c3706dedafdc5f7d031c888ec",
      x"6166deed0db12dd2ce6ecad932eaabd19d32d9c9d56580057aba5e4bf94c3cd5",
      x"a4e17a2a995e7f877d9bcf812710a8c89e174c802a16a0ef17b1980fb4e13fe4",
      x"bd0b8cef14b01fd6c016ef00fac44d0eda7ddd055387af8d5e2f332dfdb10907",
      x"739c8b2756fb6c4a38779fd9602441a9a5e7c1b46b347a3f8f3b4accfea40991",
      x"f5448a4ac9230f4379df6385bc6f0432cab4fce47fff997102f9d3da0a37402a",
      x"e3f3900b359a142fab07a4dedf72e3b5f8d95a1463861b5d9202c0536b24cf16",
      x"32c8040f859629e4d15ce7d982fe77fbdb1477384f69069b48a106c299dd99c3",
      x"fb7d89a4b9f0cd1176f13393694468623ca1dd829d75936bfd4fd28d4852d47e",
      x"9bad871b2b76cf9b50c7274de2ec9fff751b634f0c21ebb01e6bca5e4877ae0c",
      x"4fb204c12f80aa34ad9cdba9b6ebc13aaf24a536613be322c15a8b5597f75221",
      x"391faabda3d4214d905a32231207057cb2fcdf05b8561016660c2b850861e589",
      x"78cec8853cd8a5f1221edf0ccf7b0700bc6559df1865c9ee31f577da9f478cea",
      x"3ad8602ec80d368ab7b6ebb0d065e825433fde113c22a37c998b3edc8bd8783a",
      x"6aa393a896abe3b74af1b8b95670b6f724094ea4cde7c2b97bdc8b446dfdf04e",
      x"0516ebcea22d4ba7921f68d2d0eab15c48d6bfd2bc854104856007f6cda5f76e",
      x"cb22763b437da0734fed892ea91ed76555d34423c1715bd6cf8b83003f4ecaf8",
      x"ac23380f0bafa88d201f875df7d4b1a363a0ea09bf35ac4a03ac5424e263280a",
      x"ead7aa91ea1c3970152269483f690dccd188c7b911e1b16c2d07248ec86858f9",
      x"f67f78fd5518d546e16e0c39a97c33467bf22ef966aef87adffdb4852209acdc",
      x"8fbc87b571373197a60806facfadcc884d9bd34e82ebd045c117cebf59eefa0e",
      x"74cc7a76486c5edc922e52802e16820b3f1f042e1b62f1030bdf7b4a15de1dce",
      x"9faf58bd1ca44c375d80d252b048610a8ef3030a81e41514b9772b46aa0e545f",
      x"5dc00697613a32f855618d9152a660e29d2cd91ab2e90cc206e0ff65c71d5d99",
      x"ee9920a4c6dff00ad362c9c97f14c96d10485d63f24cc048ee248922e81b4308",
      x"3ad574d005c7a81a55d1f574faef971c6b82c9313ae5bbc113666b35a9e4d915",
      x"18b2ffe87d3186675513788c9ed73bc397ba20c4794785cd895de630d5d12d67",
      x"3417b94930d50525801dabf6d04c29aa0f61bd6495158500fae1ff3dbf65c5bc",
      x"6cbacb7f40c9f897adff8bb1002ccd4f6ee10978bb611480f7ec34905afab578",
      x"aa7c91e4bc837cb809f1f3ea355d3b7bd06b1bf6bc94480c0044d5626fd471fd",
      x"18d0767c9d5678d1493e1c0375daec0a4a204bf39f78374dd8d30840aa34d64e",
      x"95814523380d74e2079482e08fc471cc8184ee59b6c0dcd579f32e60bf2c4562",
      x"1883382819af8a3ef8acdda8d3245108278da6494a70cbc633ad8ec866818bb0",
      x"0b7bab69d2fae91b2e1a533bfa76e8d839a99aa74e41bbbbe978ce4a031c46ca",
      x"4aeb3ef88c2f8333e85d3e01621815b2cfc9eb8b1a5094b2b22efa5c1265df9e",
      x"f56efad0ec66941a1606f4873f977a12a78ac8cb6bc0404e53f0808980c65d61",
      x"f3c7dda0f4be08f0ae9e6d823ce236b0abacde8aacaa6945385413a49f5a27ad",
      x"3e447966b95c41c8886fdfb6b0044971d3053e9b437a1afc7fa6eff3e3e5ecc8",
      x"78bd9cfa26f86ea87f1de8a95a706f857b4292cefcaf46fec568721de9e62655",
      x"2b409dbdb18bffcd8637c0b4d4ae74d80fb2baa6aaa5b907136045aacb074699",
      x"042f734351cbd40dfdc1b406c1a7fec904a67376aad5b8ae4ccd9cf28da0b4e1",
      x"9ed9614b80da1847da8f22c0a48f21c4638de7fdfcbff128f54a23c312268da3",
      x"449076330cc37698f30aa6ca91007efda4dd0869be6453bb49a4538d9f6b0dc5",
      x"ed030d29a166c153f21232b416b94134c226b28331dc0fbab83482295ad88bb9",
      x"bfe50519ba4d82015439d3fc3490228acf70951ab41c971dbcc87b8491e81b03",
      x"741542e3865ef3a0065894d8ac1970b2e4a8f38765343d44fdeb8692c0f512bd",
      x"64fb20c50a076933f781666ab9e69fac5b6ab91afafbaa6c791d71c39a5d66b2",
      x"7c3cf9c04d0ac3c6f6bb64e9c81140f7d46851228f08e18beea3dd57d9240175",
      x"2a61ec7540f929607ff2f50f612afeb7a31db02f47208fb1f2709021f85bb160",
      x"e7c08374110fab7c3852f2e809d63ff1960f3b5f29e93b708fb0b2e658d234bd",
      x"8f358cfdb38afe1a5c7a589ab9d457e8ced277bcba6dfc770b612ae3c032e462",
      x"8ad7cf5006773ba7a4d2d542ff1b3ef9f3dd983c8c7a90cb6c9ad09aaf0d8eaa",
      x"14ddb4ac54276be9e4851b6e61c75189d15f73948b640e66a1f3de1499cbfbd1",
      x"7c9ca311e3af770ce699787381080388992e95bf2cfdb1602f2e68fbce48750c",
      x"65a395f974adff8a1a13928d7c2d566d0ff020d28ab4f537a193983a8f501a9a",
      x"3694a7ba7f234222ca12271fdd069de35f7e17121010a2fcba577cea18608bbf",
      x"321b50ffa9d458ae50c977d73245c04d57ff65973a7378ba7f672aa6e2b3e5df",
      x"2b475065d8c67b1e8b967b5fd8c391e649c5218c3b72db969aaa32431cd1a914",
      x"796beb84762903edf7a4dc054c0c8afffbb452d15e938e5ef363d79540ccc0e9",
      x"aac6511fcf252950d4c4d494d85f5cf5fc4c99ec2dccb807b859439fb7a8d218",
      x"ec7d12e61349a2a3f51b6cafb0be2a1745b08dd96358b560252ebdb4dcea2239",
      x"59fe2b7f53a720236588c1553f708e22319eaea7901051350143ad7980d9570b",
      x"90d836637ff35c289d2d761cfe6759391ab79fc5f753d0e16022b411412fc317",
      x"e2af485746ae3e13e0b654a870b945c25be789ef298fa826b9c4ef5cb3415866",
      x"ea161a7062f3cc2b6b0c1c29f5edc04ed50303a8678d8a604d29e3634a64f473",
      x"7cc69c77995c348f662b95b30145168e3e3a060914f4a79ad8b16e329d86d053",
      x"fc0e8dce0ff08b83e83ff7091e3f0fa0cdf33ce32104b4094f5ad028de1811fd",
      x"8fe9493a4b2754d72210c471b9fb83b4db4611030015889757a5c86c3cc32068",
      x"08127c3803c08dffbfd2162e84033887c7948ece34f6b0512dbe262d608ba194",
      x"a6a9c1c05f38adde232f2ade3df65f9576404354a583c3828887021f8c5a7459",
      x"a2f402d6249338766533699f5a6196f27b9c50a4443c9a960a429ce51e2a2d63",
      x"adb1fce2ba5658db6b2404a07f33935b36d17cc3f42f23a2a223d40b5b229c10",
      x"08db8d1bd032300a0ad37839ca0c3ddea8c4276fc08a4970a1b5878fffef6a9e",
      x"be569f846d9108420ed3d7b12a9021782b2aa57931efce02bc9097e5afade4ec",
      x"d6e833bae8512ba5513620d3ac78c23b6dc8a2fc4092ee386d0c9bc4e547632b",
      x"7a4cba8ff195efccf818c7a0529084b9a1beab387920f1d47489549cb4426be4",
      x"00c0a71cb7fb3d711d9298c91440f212f8318caa925f96576a7c47ad4eeb7252",
      x"825b0b0a41b84911072c040a53d6bd8a7644b11bc4eb4052ff9b814e20f6467f",
      x"8d13e7bd4c8a31b65b42074f1a9ee2a468875cdc02025741764a092142590a17",
      x"fbff251d72a22c1287f0c115e801c3148490acd0ac7492c42bf0af38d3bd925d",
      x"f6070e808d7d53c41e14889aac1cb251f831545e83e64ee855e70ebe7057f0f3",
      x"bc44fe8dfebb3c424c65ca264f2531010a5e1caf44f13d00bab0d1e199f6ed1d",
      x"5784f1ae913d55f3d3d2840ab050faaacc83fcb4797e7764ea8b38dad4f3df25",
      x"69bbc89f038296e2ee2e87a3f00aca6cb01c70ec05a934201223bed8ec1f46f6",
      x"0226ffd47c1d29699d29a8ac34c30e0261f7e4d7c10a6ab1db0f2c94091329cc",
      x"37ba61ffa5f673a00a00fc8aa3869287dc559b34d187aa35eba6321cac1eaeac",
      x"e051ff69016963f815bd9ff5546cd66ccadd98d0825f5a4881c1804e24bf28ef",
      x"84244e908e3e45caafd4c3323682647a41e2bc7e733a5716a6de337be5033fdd",
      x"69fdc95c605b2b7184e51bf77452e01481cb4068fac794f0b096db41204e0f86",
      x"fafa2b704d6eb698042fb4051229063d88b8541ae902d54bc1508f88ddccbd76"
    ),
    (
      x"bbd277df4800ca1392c74023ff95f33d55a6526e4c54046b0bdcb3ebaf4e4711",
      x"6e82c88cc2e05fbdb46d2fa69ffb698c4afbdf9d9b14ce100273507541cfa561",
      x"ba9d5de75847199ef738d81fbc3afb9fd7b38a6d46ad0bf30115cefc7888f897",
      x"f70bd1423edc066dda5d51d665a24d7dc8760d5e19e8375ec8dfb1b556d01573",
      x"a31b737b60e79b129a3a8448384afecd9991a0a1a226f61bad5fb2755661b9df",
      x"8fd84e19a7c376939d5833252070e1801754f61fb5397c0272b2e92c6bcfa7fa",
      x"00edaed933258c442924d8bba31ac4b1de2b9fc5ba926b82debf4fa28f1d2ce5",
      x"4af113bb82bef6d8e63f161a0dbd597f1429289bc841eb73da8a869ee1286049",
      x"3cb8244faf976fa0db879883ba73e376a3ae08867e79b4f7e7b1e9fa0e8f72f1",
      x"5cd9bd754d5fa758d431e0e22f991473f358895176d7c88ac46535fcae4bc778",
      x"e1dcd9003cf4fca825ce0f0056beb6a0fb0d1a036c9e4f0d0e624fcabb2372e7",
      x"76b1366fd91cd2aa3af35c2508677716b3b9134c92ef18049dc786a74e4ff9a5",
      x"f405e12312b0f73ede59427bb8f8bbdf026d8573c5f6f4b909f444e51b6f3223",
      x"e637b6abeec2431f2303390252cd03f6d30ba1f49a40cd6700736450a03347d8",
      x"7587141e76dbffc4388fdb19e34d29f34f819e220dd3c9b470955262f68349ca",
      x"e3b5c1107be3e920f3a87067e51ebdaaec9308f230fa4494e2e18bcbe5ffb2f2",
      x"db7bda782229f6296ba706280dfbfbe6f542949802f66cc42826c74169352860",
      x"6b762f59586d642a49768662575c9e35ea71dd5f7bf503a64e9d62b0f4709fe9",
      x"0323c912a2768b47eea91392de79634cb754ed79f75b3dc39ad9399723d5a4d1",
      x"c4e8fbb3253ef084d6028b2c27fbf07f332a50395904b0e0e6b36cb9623faddf",
      x"ad83fdb45f400e0d8eae7cd348b6c69314476c05fc6d77f282da0df472145adb",
      x"6c1981bcf571560b0a2583ab1040085a753b13a8b90a17f18839ecee5d179bf4",
      x"c08b22e5ea073286416d69d03095d52f3652ba0d2442645b18dc5ad734a18c36",
      x"66808c7ee6bf8364f6f2fd819f59d2782ff463ea00babb669db6837ecf4a7f4f",
      x"fe627df4f89e9eaa4faad8729b5d594d1a5cfb42731dd701d3fcc01ffed8b0bb",
      x"82ca211059a6940e6ddcb76872dea2bbd1947fe9b9355333958fdd0dad8765ad",
      x"4a99a5c9935d46df23daaf97d80a3b32c5f726b253b63b02ef51540b0ec04ccb",
      x"ca6d64eb3afbb5c11f9c6f8f2e90508d09fe9726634f669a93d3049931ae5827",
      x"7d860c38dc22a06cd39ea75a90b22ca2a9fd870dc31fce3b9e5c61bbb4a698da",
      x"c6b4b60a7c8acf157e890953767bb97cad0a83dcb3a8761bf42ab57edbbc5de0",
      x"09bbc5ba1ac0bb83ade5a94f75f578b17b0106b25daa9302d90c4e8439a02edf",
      x"3b3268eddaccf3251bffd412671723ed056fbfb9fb06d989e176673986a3629c",
      x"c9407f491d8380fb232a6827a0d2ae53e81ae08d5796a1288790a09c0e5342de",
      x"1fb3a755901486180125b1219fbc20fe7232c68ee969af1c59f296e47fd63112",
      x"8cd676baa9cb6e9f292ebc34d97bc9cd567303cb9bd15b9fe036e917e394c6e2",
      x"b0f14b1bdb7a11b652aa6cd56c6be04d2866db38c043a8ce7aa8bb43b29d59b9",
      x"ae0cdb86bf6664ecae906fd9b0d57412daeaf3d528b61fd468daa73f660ca38d",
      x"69ba18b95455d9bd09e6dbd2c966d61aaa22dcb6f6aad7cb8255f657634bdd4a",
      x"655869389c14555b9d1b340b67b2a078245d875a873cf4de49e318df5c89540b",
      x"04161d1147c51abaf192c85f10acbf91bc1fa363b9bb5571e632acda1efd6762",
      x"8e10d75b4c2f6fa3dbe85d9619d164b20231c25250e3dd582ae0d769cf9249b7",
      x"957ccb018aa92649739f4fb5a0cb2bd57a5f740103c7be5fd3ade3cecea5d4cc",
      x"449ab37e3438924f8f0c2af511a45e6ea3776016b50cb3d60b6c981855e4af83",
      x"00dc5a3de57ecabe4a2117657e70c98a98763d0bf83ee09a01d60879ebe460cc",
      x"5136c12a26b484c9212430688b53495c7b87090ee7f520908536236f90d0cca0",
      x"c4460c262bf78e8e5dde1e38a63ea8c443991e3b1fa4497ea1dcf02eb3c935a0",
      x"03af2a7fd91471157040d68db1c465f9c4a0dd475cbe37ff23bc35a0db721ead",
      x"b1e539be582b999e91dfe2db179102fac4540739d56c4da99fdfc5d8b603a880",
      x"f579063337330b8e3705057df55af3f804cadd674feb14d3008f07716297b822",
      x"f47c73d0a81ecea1ed8c7181cc2a3650f1b362a630e54b42bc64cf2cec9b131a",
      x"f3287a9e2cce248e71f7a09ae8006f38b41fc0da339f3c6e77eb989ca2c3a49a",
      x"3a8a760d8addda1e2a343fd2a5d505e9d3a7e23a3b8628c0c8f632b4c9a7f2f0",
      x"52150f05db9dce2b22d8fbe7f9f9c345459c9cb7767d8ffd73f2898dcd78f7ce",
      x"7f7050ec36591685923f40bcd8757a9097d65cb4728811d29e9436190720bdbe",
      x"86cc37ef5cfd00cfcd8174d779451a674a8ac6a0aa5fafe49816fe778e0bf2ca",
      x"d8ccb84fb9e331252d5e9d6c604021cfd6ecc46c62bbcdf798d08240d7add77a",
      x"9f948089290722b071983cd4f63b968a3cffaed800c8588a46f4d7fd2d58c33e",
      x"034bd23a957cefeaccadbefec6d67b3cc943906828d86e5693686d144740d66b",
      x"070d62cd533e76738fd089690b70786ff24d799d9a72b01867a5828831ada629",
      x"dbb2380070b15f25e5786be53d4f983ab4f2d5105a184c917bf4d626e7b68465",
      x"c8a3f19e98eda7368a13806ccda32d5f8817a2263d07537ebd5b0062133335e8",
      x"93a2116dcb2bed475c8cbae27f89b0835b3b5280c040d6a9be4ac9d3411b9f5c",
      x"6cbef64eca8f04b8aa672ddb04303c6c4bfe0b68fbffef8e9685429b4a09b5e6",
      x"103ab3b21830cd331af607ff3ce16ccd60675d29a5b6682aa6747b5b8462ebfd",
      x"b4575f0ea0308b59c723945180131caf181f46487a9801868de6007a02b5ee0e",
      x"a1bf044b70ebcaccc5f9de0c7e90baa834c9f57e6cf3ba01b3a24c315b5fe360",
      x"9092afc54dca53b9b8bc694f12b44bde7ce09d60a86957543fb7f76e95bac9cb",
      x"d3a9b31f3462d9acfde42db30a4856c43f95ba8bf0fa5fe8d6c2cc699caea3ed",
      x"f62f11a3f7d6be724298de3c46a02040007db2126406874f25bf80d06f65aae9",
      x"113c2ad5459f2ca04b9c82aab8133528e56de784d0968ea45e148dcc19bc5579",
      x"42a60d1e03c4777fc1a3a75f302563ce808c5ddfad9fa1a2491a5660409608d2",
      x"b05cec76f9794a6349e74d456e44789c7849957b8d3af9b489e620505c69b835",
      x"01887843d4c02fa76823d65dc4ea5ba4478615ed9a01f5f64158a7f0b683c943",
      x"6ebcbe8907683ef8425c8509228fa5df804a7458c043e64d33bb94035bf9db47",
      x"5d9c4f3d3558b9a531f013e05f91b017c35ee2f2f8008d2f05e44a1410ef30b8",
      x"93ab933a28239de618b40af4e6b961a80e8cb369d7398b7723c8a01e3b8d2fd2",
      x"8217f3b8f27f6ac7fae7f6403cdc769b4830137567209167fbccf72022a64b08",
      x"05afc3966bcdb6ca1cab6d8f6fcdd474256fa91f8686edccee23d652fbb8464d",
      x"2353b256da7733019fb1cacdf67ad46295b10563a69c15c7bbff839cc1590140",
      x"040287a46b32be13161a085d5a4f88c9845f8b351bea671f1656222ddc01a094",
      x"ff5a3242ba81b8f632df04c7f72e0a00b9ac48fb5e3f5008ecdf6ab8ff958c38",
      x"32b60e283f6338baaace6fe1a4c8806e1c0642a4006b3812dc27b24ced099575",
      x"0e28ec98e0d71674b959b7ccbb29a12edf87607549297b3de9f5df05230f3ca3",
      x"0ea9298fc8e1dd30c2cfd6d872423feb16831a36acabefe59d3f31bf20537f2d",
      x"238c97eb120a936a5a8f835f66cf3b60c0b7f33d8a735bd788ddc74f85c19b77",
      x"7b182012ef6f47c2d4cc8bf31970146d315eba2d132982692daa842dcdef744a",
      x"5b96001b631d6d14c7c2e843c03954f566cb4681ab3072005bd167639fb4eeac",
      x"08a6b91b6c3fbae4286f9d2e99085397b8a9a85001478d911a3f2620a1c22fe1",
      x"5afa335825c60d2e87f57f9439a393de6d604b37219e09f8a6f2825151cff810",
      x"4083bb6771de955dad397a204486f478df1be10b7a288efa93dc692163b62ddc",
      x"44ddef11a246d8467b581a18717a5d00b489cb3c61ecd7382bdfc768da7a47a7",
      x"5ca7e4624a6b70a0fc8840a4b453e0beb0c7f237c1b5ee7301e4760257a7ba1b",
      x"ecfd259188ccf84658006c8b98c1d56a6daac2b4a8caa35e8b453cd2d129c9ff",
      x"a0252da7811ea6c908bdd234d7bffb900de84632ab4e5c78f04c08dd1d93b982",
      x"7b7b9f44c3678e7abbe8d7520dd018ca9b043a993a5ba964fb7b7b678e1d8013",
      x"5bbb0d5e3639af8025784e5cf5251ef5c03877bae8a357fe5b2a8959b8ce809c",
      x"7a9e797256ab275f93739ce4038a16f9b99f5cc0bb15c9ced4f93722b94b91a8",
      x"70f752d200af14acb1f10fbfa6a2854a8c10c8f724f966dfd4a067e9018e3273",
      x"a3904cc9904dcb457151e56e4becfc04ef1172b68040de240aba0254b9e598ed",
      x"fca1724cf0c32c36ec75a4431934b5d4e5248d2636b5271cf5da5e996b01e089",
      x"253fc778b5e38321f38d4d8f91917affbc9d070e41e0058f0af176a32f87b899",
      x"590dbe7a3fe7e5d800bd3381a37d62483b127feb47e0545624ebceae0d9f27b5",
      x"620867f1e1ee9e2682c5f6b939216aa6068ca7c93978fd5a736c966ac247b80b",
      x"f98d5ece089b6b7315564c9e2136871ba489bed231e8c6922a09a1d170b784a2",
      x"8286069d1502ad40e37270b2b6e3c30d5c13ade819b2650652641ec1e8e037f8",
      x"5e5330a34c1bec8fc4974ec2dc85bff9f97b4532a629b822dffa25e261affb28",
      x"b618a7112eb1360dc39c1225dd05b32c8a288f4f4b2e60cbaea7129ca8b77782",
      x"17dbd27bd9637aa0ff556d4c66ff27d8c0812fca9eb6611525a36a3b6598833f",
      x"f1f75450fb8ac240e1f985ade2c832edab241b28a95afad13c4f1af668c0155a",
      x"b1e6a630d18357c55200e83347c350f1ea31e8935723c642c2dca645b21a9d47",
      x"e152e507e16abc4d6a97aa50e21cee040b21518510ef8ff7c37de06eb218400d",
      x"658e6e8c5ed0732b66d8a89e98e2890ba8800abb54cf911f227fd8ca3ac3e3fc",
      x"23d7cf21563acf539e42b0014b19fb2c39375e36edaf64003667b6f124cf00c2",
      x"11acd1273fb416fb5ad3bd8227773700a0d2a2e15545ea4d58ede2d303a6925b",
      x"bd5ba88397794215bfde93a30d9e3c28512abdfb9683200e8e9559538b5df08a",
      x"a822abb27da5c701dce0d8592139c08a7a9534ada196a950ee413b3901d23986",
      x"51de1b6f54de115412377a3527db13b399565f758d62ede9007dbbdffc6c787c",
      x"b00edf1f5565d3fcd76ca15184be24cb4701a03568aaf464499d30744b1b83f9",
      x"259c7a25bdbad809067a4b429534ab864d959eec55faf41a73c698796190f531",
      x"78e4d5a131d2cb48fb9fd3d10236e6695812586d2368bdde1b781ad43d4f2c93",
      x"5560b92364ce03e5e5b8c799685da9352cc0a0b0881f4a676634be4cf0591de1",
      x"a1ffe7bccc8e25c634a6d2333547949aa28c756fd9b610f14b8a76d2cc221d80",
      x"a7fcd9210bd38a4bc7399b267e54af03ab021aec07a9164239bdd9f0117137f6",
      x"04513fc41549da455b66ba6646bc4075a07d3cef86200f7f15b36d15a42e49d2",
      x"3f5ddeffb581d0cab5c7f77bcbec299d968ef48576c82ed3ddcf46780dec23c5",
      x"fa353d138e23c40b5657551cbf0d7cf668b34b40a74ace58f868e94f7daf9314",
      x"6451cc3abac26d41e8c600dcdd821584123444e1b478126272587d93fc831f67",
      x"c81d55c0f6b0188ca878555513b38af41c26401bd92cbfa9060b38ee5ddbfebb",
      x"1b4c1d5fc0f62ca29f7c848b131310f002f0eb0db9377523203c4200724e3f47",
      x"736ba32ea31bb113b51c64d6f2fb6ed40dcf9b4bda0eccc588ce435296d5b3fb",
      x"8537a95d565ce95be1c0757bdabeeeab11bfaac13f60d224137c7ee292766b95",
      x"aa1b4ff5a7bd1e4787410902e1eb9df8bf3c7e76805e5e0ae8ecda95f4f9e2af",
      x"d9931dba44724cf77f2a971003e74dd447278ad9d489b1afeaa20d3b026b2c2d",
      x"37478679132e0f61798e45d95e9e49126c3e9edda1a469d607f8d6d0696a2990",
      x"cd0764d1867bc82feec4f9717d090bc710ddc37a319d95411d01bc19a4cedd95",
      x"3497e7197ed45846fb5edfb2409b2a98817904a6244bade231553274ba25be8c",
      x"ec2427e9300425bb5de6d0ee151d74eb6a5ade25bddbb9397022a5344a6d37ab",
      x"99cbd4d0233d295aa743ce8c6de96662d8d5fb33bb5f34e550f4495f0f006adc",
      x"1fbaf6bf2623c2447e895a6a3eaf12bec5d0716c85fc2759d1c8b66b0021bf67",
      x"48b5f44de00547723417ab1b15107dd8b12bca012b8e756ced5f589831683ceb",
      x"059eda049fd17c1f44895172bd8274cb2211142648f22949c77357fc2a34a190",
      x"68619e93c7853c27027abbacfac22c26858e4f3745e8d5dede7c72f5ef512b12",
      x"21a254a37c4f1fc2cb639098d9fb32faa2407eb8f9b2d72930749fb723c5006e",
      x"ce1811da26a2292ff496789d4f84dbf733984ff4451ae2cd81799b4d15178a01",
      x"ae52e2e5e9e551f7b4065930313052e3432c6d8a97c3fca05e88b576dfe8ee96",
      x"5a73c849da9104cd2ea5ee065c2389d4e3fc3fcea6a9a3d904572f8e03e62c4a",
      x"074b2142ea2bf78eb40e0e86a5561c956c18eb8edeab91258e5507d1c1b86afe",
      x"49b180998ed5c436b8297a6c79325edfc3b13fc939be164f15f5ae2b19a4a307",
      x"6abdab1a1ade24a95aa63dba92a9d99a5f5a60dd002c81d90297267c96159424",
      x"ef9c23ad996949ab132739ac32069e4b0a38518cb6194cbe1ec4bedbbf1758a6",
      x"8c12388c19fa61f3e03ec24b438ea1b3f114144171947310d2a965372f5ca322",
      x"77a1d061450333471fad08a0955490d0df6567d78bb68e094a08a662c46c94de",
      x"a0ee81086b89d5292f13dc0f91a39ea15bfbbf3157ab0f55c1ebda010cba7aa4",
      x"e070c9e788715068b378edf25982e1f7158a08285cab26c2ff54007945ac8916",
      x"573da046870778d58511272c145e0c2b349c5033ed655cc5c92c82c8ff9a42f2",
      x"b6d160c2a15eb0db3e2a565277ae8129f6516f0f98fc8c027c607c61fb05a844",
      x"ba479425f9ead056da987fe81a945b77e1e695e2b0bd2b94ff2bc8c4b58efeed",
      x"734b083fb53584625a01d099588b64464f50610f92f7755ce2cc666a1bc1720f",
      x"cfa56e1b8a3d41fb160d3ddd660db7e5eee31e94998ebd591d2600689d566c37",
      x"f37e154c12d66a8aeff001822c2ed294f54ec64832426608b031c2e9849f4910",
      x"d054b7a66e92d520407e3eb27428789c645a69b0ffdefbc0bd106fa52bf8406b",
      x"6566599300ddf40bee267674371c78a4cb3ea14cd44871c20d9410b5f25ec8ff",
      x"9795fecd5a63880fc289ffe0f5a6de8e36880bbf7568c92fb041d934491898cc",
      x"1625d03497e53b4ebcbc16757139cd5cf620fe7b61fb366d2429f58a2c42946d",
      x"ddf0f474856677764d6a2cff0d92016da60845385318265038edce00c2ebee8d",
      x"087eb16a9f3baad00f878ff79500b9ca7be04829ead02e8ce50cfc5bb7d82b8f",
      x"531313804d27d56e144815832cad01904227b132d4da4b7ffb63e1a2e6deb7c5",
      x"81b51a953db853f3cbe342ed6232037d87776d10762c78a3f3ee74755395ab98",
      x"8d2260e15c39ffa9ba02636c3589d18d479558a81546fed95f4b7df10a74dbe7",
      x"f0fb9e632f63c3aabdaf83e812cbac69b9e5bc737b8e9cc979180ea0836bf624",
      x"64cd84fc0db278997eed6d48c51adf257227e87ec89b34cae2e95ffe0b55996d",
      x"170e0cb3e109672526fe9d0fdabe87dddfd8dc3f3df50de2bfd108074f1f1b1e",
      x"40f76507f96eea722015857881da80f65b44bddd27936284af8ac277ff8ed440",
      x"f556abc9bc478a510383df105bfd150cff18779c76802c292282686cfb6e1bd7",
      x"b64c2bd8b47f184954681aa830199ed05ed133c78db52d270ab3c22c897c3c3c",
      x"346073e7595320ebadf6ad749541fadb4387bf8cd5745a90a7bb6797ad3eeb2f",
      x"ca091320ed0b2636087c132ec4e21901c66adb3543613738349aff2c37cc9d84",
      x"7ebdffa3e997d39bc1ee8d84b84bdf0ed311db4c3078473436c3d2c9ff2bd3ca",
      x"86c6aa68be91cc2ae6c0c2db57203b5d44d07681d77d9aac288fc37f19c5d9b2",
      x"9151df1ff910e49db5032b18452642ea31e01d457c22e3ca609549bd70efb828",
      x"dc5bc975d6f80add3d74f36e719085ab391a937f8c4abff9b36c42645738fd8f",
      x"5cac9decd3703f232e4e3757793a290530821e2919415e6848e06c19f1980b65",
      x"dafd8c96055e5c7e4ad1cdc49438e246849df1a682baf5dd7e8dcffc783d26c1",
      x"22e3934fbc61fb22ec9e87361eaeb89aec5f423c8de7cfaf70059de5d536c6aa",
      x"b8b7b40e0b6869393d1d4f5d661d6bf87ae4b35439cc1ddb10b7e94cd5ad4726",
      x"15c50f355e3d2e58d8c853a29067cd342a8158e3f2c0bedcae2504f088a1519f",
      x"26882969e5d5918c48651c73cc46084884943fd4293056070e192edbb7b8a71f",
      x"0051fa809badc69f7845d1ec6744787710b00effba2a149795dde423c8ce1df3",
      x"e4a6b4f558cc7b79b06494c9ceea5600905cfc93a24c0735eb8a9e64edae9b39",
      x"a4f29f8308915662a6ac68b2f1f589df8281620a6ec277d58a6a78e7c2fb5306",
      x"c891114b93d4a5988441289abbf86688a841f87ae02c2501d1a82ff0cadcd9aa",
      x"032f81d1fb7f91e3bd91b13e2805b757f031ce6552ad8f0e3731a100a2af2f20",
      x"fa90a53d6be913d76827ab8accc0747fae4ea1ac0b7397006d24c47ccbbba0e4",
      x"a618bcaedf312a8e11e3f5ef4c3a072a11d4afe1f9b360997bce94a870f234a2",
      x"20e5b7cb5096ec430b28dac40aab0829b25abbd2b1b2a146a4f59d74b4c8097e",
      x"d64d559646b71bc9caaa0dd7e2f50858c580572240d703d5bbeab4de74e028cb",
      x"f6c6fb8e73d9c00565a473b87d10570f373d5e1638fd6ff6819d542d241b72a3",
      x"738ee63e3db41e2c7f4e6f85fe50a52d1ea97be12d0b77860b4183bb2bf60f46",
      x"61e1f23931dadec574962b7d3bb9a6b504550039f785f171e95faf1676303c59",
      x"62aa039c03ae76507d05ca27d191974ce1d3c951a414217e1e1c8c40eca22168",
      x"7399e86d2641626a28981ffbe70ec213a8523e73a35b930fe04679643be2d209",
      x"7d755875b7185570de318ad37831264bddb2a352823b624183558f39d07077fd",
      x"6f0e861dfa65d0dcb4814a5f78894b7b2ba0929acf2b4d1c3b63b9a5da65e45c",
      x"52f55a1695011c447ec90cb9c1144ad52b760ac77aa8e43675a185052e7b628a",
      x"0e8a1c132fc170988d404e8ac69c8162524ed30d4962bdaa89b827fd3fac514e",
      x"c6163b97b89d8e18478f75e3b2ea1255fabf4cf7741e81a452308899dafd195c",
      x"0cf377dd58dccbe19b514dfe35d0ee168ac86eb5591e50992d34b97f78fc327a",
      x"3b722ef9e6f17b87dae545a67b40230e6d4e24378cbc5aa33b10c1315e6cde6f",
      x"0deb3e23a29b8563ac4933b43429c7016238564479bcd100ed94ecb32952d4ac",
      x"ebb69075b3b8850102da704b9219257f1a8dc5a811a8801148a5b83071a42ea1",
      x"8c47a0e255dfed03a9896544a2fdee5ce9cc8ca9b35075876dd4924738195196",
      x"c6e1a0b8c9d74e155a84f43fc21d61e537a74623cc5e3810405bf2e86e4d1e3e",
      x"0930b5fadabb82f8f9def282ee2e49351615fcba2167c6e1a61663db4df55674",
      x"422d0a6de9827cee6678f70d86884bfc4c62ab53fa644b0b076507532021ed91",
      x"4c74d0a86d3bde9aff9f1c27db130149baa404872ccafc0e4895d7cce300ce41",
      x"4710ab966450966e003bdd5733cbc384877e4daa8f706ad619eecb55fa42a039",
      x"2cddb3834dee4f5a08fdcd05d404723f2d1827c9ae02311878267ab9989831e5",
      x"0ba1c292d964da36a78bf54c6d59cdec2559f3ddecf879d95ab51642ce61e6fe",
      x"5320a3c75e161df56be3ed0f01b7b18dbe4eaa317b21ea507d98f9dd4885faa5",
      x"5e23561bd0457ace8da62fc929520de620d098d945e780823b6df4d3173c5abf",
      x"9558b533df5a57b3eb5b3ff0d831436f5fd4a469e87ee952afe1f7f27f0cd2aa",
      x"db0b9429be911b9de6ee9d5b183e146dedfa3c435c5a740b6fd17248b5b0977f",
      x"ece7b995ae836c75f4d484431099476e7da1c3133e829422cb8363b1337538d0",
      x"4f3590b6ff80562674212636f12c99a9465fec6a0fd424b8494140c76c188abb",
      x"3a9322a082ac77742f21d60d667fc272a8f3ec0baccf2c3fa42f982723679a51",
      x"3a7a7da533da826a5a6dee9e76d4f4dd6ab44c9c6b00c27bc7e553c2fb8e4948",
      x"1c605d62b3d27545d5e59d4554141dc889a952815bfba9320feeb21644ce287c",
      x"cd1d81394558a048fd02e9234bdb95eda15b0156b78e64b5e3170dc09333e48e",
      x"2d32b5b11e65e0db185b56cfc01bfffb436dda3b5232ae65df5c1ed7c5e58a8f",
      x"8d93a9c8df33fbefabf14616d3933f38c573fa0b4ef702c72ca0979753aa1bb2",
      x"db304dc0b6886f3f7730e0436e7c48de7c825baf58f05880a660bcc6b9dedf21",
      x"a93ccbaea4b59736977982db82497251b80b44ec01b2961ff74d61873a262f8a",
      x"961f0ae8c924326c47109a5dcf0f92afca9ce7127cb81aa8e67a5021a86247da",
      x"620568e81b28421fe379453b62bf6e7127eab5de3a3f55a974bfe70e0f6186e6",
      x"4fbb0c0d66280481f21223e79075e883bc2e4b01db7b76841843d877b12eb556",
      x"02bd94e27355a0d42c740b83ce71f37deaffb5c3b61e7aae6d8eeb5045fa6d7d",
      x"98ce952de1f78bd1ddcf1a625fa8537c93661a9f1121c98ea582ab2f99408551",
      x"80e660342349544cf0418c3c266b7578483a8bc3fb6906d9386e262c14d72a28",
      x"7ed4e6df3b51fd64cc1b87fdcddbd28cef7de6461c6502de0f26c89215399e7f",
      x"df48fa83eb3799de114dcfbea09c33701d9aa57e4090759370e95830fd60b8a7",
      x"d15b1579752b50c2521233c2c6e214afaee1c61ada7bdf07757adc6bbf9ad323",
      x"13cb3d57f87667fda04370075002aff2a1dfdf48ff1af590828ac494e78bb999",
      x"ce9f5d0380ae6db07166ad3f52ee8dec3cdc91f558aaa8efa74b2e023fd39c6b",
      x"7dc86edb8a4fe453eefd0b5e79c3e2efb05050e78384d24f61f273e64acf583c",
      x"1d8f11485ae4137911a60bc27c89219917bb72e66ae2bdf2f2915c6383790e1a",
      x"6f4a1c3437c6b3f82f97da04c71daed01846dc7db87ec7d2ccb27d0a9fd2d0b6",
      x"9b3971dec5b3ee490bd807ced6d1ee74c49f25249d43b4b1b01e39666a340d84",
      x"554d6fcab9bc053ac35060ada9b788d0474e3dcc8dc52691067706c43e2db95a",
      x"7a50ebd516b1ab676c34b4e04e44e8a39a9dfdddb73258df740c772074a1593b",
      x"ac2cbdd1130676fbaae0faf180cadd98da4b82e9ed0a34063a7c66f0553abd3c",
      x"30a560d8166754e2ec6dec1fc11e60f8c43045d6e5acdf309c9613de1b8e854a",
      x"5059c60a79a62936c0f5be04d01ebfc807bb84c1eb1e8b4a3e0e1841aa5a7296",
      x"bb6aa72ffa7245c2c9b38e64adb502f1d2fa0a0c999e938e6675f6c6cf78efdf",
      x"2c0894fdbebf270e0c332550ffc994309d650049243d798069013b5f965b9c40",
      x"cf439fdb6a15f0ea01625570e4ebd4b9e818db0ce68244180586d93c5aa3a575",
      x"7a557e1d3a9b694b7d6ebf40cd241c9ce12bbe30283134baeb7df36b658c58b9"
    ),
    (
      x"c723bd7dec784f8dba0b937c571801e9cc59afe2258f95d149600d15eccf375b",
      x"41a2feebef828bf3a9608df09f9b8907f8f6588f4c2e8827e972992718d30529",
      x"ad0b9f996f688c3729e981e53fe5aeb48ec9e5220afb6e6dd457090ab0bc8145",
      x"e525bc2452a6fd57ccceacec83685fa8ae8994d5507ac4958276ca60b515ac28",
      x"c6a7c6829113915092b3678606ef2b774b0fb0a94320bd2243aac431cb13d90e",
      x"6a79ea7d26691b5771e646eb845def5cc567c4fe59a71db3639a47dd6c6d0dac",
      x"fa1da919efeaf2fe2012dbd14ed0b5511497368467f975cefda094ae950965e1",
      x"e8cfde0dd83fea70d20fa2dcc290ae1cdd23642bb043a6f936cff7d05da8762b",
      x"a6e1b967ce4e55269e89caea404697244cf411fcfd3492964234ac27dd3c2be5",
      x"8e478e3c1787496249d2602acd1e5d594eae17b55f68e129c4be8b0aabd4c3ca",
      x"18332e3fcc9f2821345693d5394d62197a14bcddf52809c77fb40d4352683fd3",
      x"4ba5154b74dbf14c30e75bd36f0a1f7dec0ec4c87ac654b2edd53c24382dd75a",
      x"52fea5d292075f99efc6586c620e83427935678f019a218756f28ed8b98e0889",
      x"b7376255dadebee3c24c22179365161edcd1159f5442d4823b011ee183af7687",
      x"43ba37abc96ffb25cdc40180ccecf6d711ad52ca5798ab5d009c7825ce55f23b",
      x"d9c65c7f27692833d1069f6910ee9385ed1843fe09a4b64f2afb7a310f9553ed",
      x"4a0ca35ed2b3f4d926e4c905129a6e29b3c640bc51ffbfe35628595f77b5702d",
      x"f19a4abfbb13f689adc9775ecd1b6a47fdcf4cba9b4f72439ad071fcfe29aeeb",
      x"a8d11301fe6ac7d7d1fc5437138137563a5a9a0dcff89c595768f37f5506a685",
      x"bbe97b03c2cdfc31a85cf405147fb6720ef4489d2bb7c6061351b41d1391da03",
      x"1cc2e67457345a8b68e307a498698a8d18d8cff126b174c0918a8c0d7df60a42",
      x"ee41ceec8c48332d9636e0f52365bd7d15677f6dfd7a9838531c9abcdf7ce360",
      x"3743d006e4a1e816b1254c0741eb673ef14d5a6a5e354d91c67cee9524369b45",
      x"05ac2afa6e0e9909eeb2cad41ee63f50efc96164b7494b4ad0c610e0c51db3f0",
      x"54339c9edc43f51cc1a485b94139a792cd3deedf0deb36aaf0a760a6cba5373f",
      x"a147c5f245ee83c540e1d605bd032c6caea1e3c724312b5358c5a14284f4d16c",
      x"ea2c3b6a8c27832a4e45b188a047844bfbcca876d00abe554257687313932a19",
      x"84681ad0c649e6c870ee20bccb9c7cb03051787f4362011b3b8c412b217e5899",
      x"2a539d3146644b11ba06d1e40f17e77f8adc9624a06456e2580063f41bd2ea4b",
      x"903e13a91e0f97fca09fae03a75d34b47ef264633b04111822a292158fbcb6e8",
      x"36776b66d464ad9bab8764373604ba5dd4622c5bfcd29d30be277343207fda11",
      x"3ba98b1367dfb78d7ac182e64de09795ed52684fc5bd134085de967634651769",
      x"3da186f309f9ef22c4575cc30a633ebcd7e60a8485ec4f5f09e1dd108efa349a",
      x"09bcfc369f52d250b2fc2ded6daf5ab2f84aa58e978ed3b86d573349ee106e69",
      x"a37fda837030a8ab44fd5c109b04fc134f308b2f72a333af467e0d54b7e42628",
      x"9a8ac7f691abf4f6f8e3c995661fac3820373ce8cc4adc8940956b19ff7b1f16",
      x"bcafd78d0a9ea25a737acbdc1117873632177be0172c4699c6617a9e2932fbdf",
      x"6f4bf820d73f7235c371d8637c81129e992ad3428976bce94fdfd9b11d97b01d",
      x"ffd760c1f7fc556b631f686fd241d40d77936bff31c3ae3f1fa1d80f661e924e",
      x"85f6c35c79d08a444cdfd315be940b6984bc792656b2e90afa31697ca1e502c5",
      x"904c286f0c97607637e8080ef1e957392ac861fd58455f64ca386b1a2df07400",
      x"115875130fc24a4b5650a5d392fcc0526c62492826070f24ffe7bc146c88ad3f",
      x"edb38631cf641dae93df9d3e242a90c9d5723646468b26e9751cb190fffa37b7",
      x"64d965b9516845bb4ce3a0f46f9400c182fb9e3c0e1c678711b7f96859f922a9",
      x"327ce4ff4707481c734f5459169fe2ff195bbd94efccc00182526258a69268a7",
      x"3b6d8f048f5393f448e0731725e830f9b28ee8125a0a1145c21147e118a8434c",
      x"d21843b1290af35ff5e041ff45ad3ffc03f2c530cfcb44fdf9164ddde4039daa",
      x"24b931eb9ad66ee2c68548e0aaa468ecee888f002e748294364f9a0803d1147f",
      x"94661c81635d79c2154b6451f3e5427d0524bca0777fbb245b40febe174ba44b",
      x"06d160467984655ad320d215a5df1e012d764dc82f03357b68bb2ee8e5f3dc4e",
      x"0a8c166a00df67134daa2b197685040f5ba0dad69864a6f9c83072e7bb4df81e",
      x"d37e092cfce0fd11c53a007b82ba335b6d4d524c06eb4c58419f85a084e3da42",
      x"1def1888a34159a39f3404977c58502baad8e9d290c6a4547b0cbd2bb97a6b7b",
      x"90006d6b9e31de7b319bdb52f5e18ecd4a6de46bbd3c95a704feb2dac496eebb",
      x"c2e3fb24e574c6f8c8388d5e79f18872aca72645bf01df0456c1db9ac375e281",
      x"86f676b970b1a8339e0a1f9ee35c64106b69232ca66753b5bf33f460a8b0a93e",
      x"2387b75b96763b197a8b24eca8c0938214185a256e9cbf35c7b630e4d84e678f",
      x"4200052ac933cfd033cf83d8447a079c6a9862f89d20f40f592def5f1f86de22",
      x"bfc48a4d21b6f21259a5f9b42b0cf842bed8544714a59bd662647586205e8292",
      x"bf2a6557aefd6859b43a33868c64c965347e6018c699651fb5a40806f74b0398",
      x"2e00d3cfaafdcc440847e7ee7fa4108f77195d29184e3e3aa1a00a0a373f505b",
      x"168591dd627c0e16990abcbd8e81711bfca44717659c2a642278b385df769002",
      x"52b9564c078b673afcf0e5dbc86744e97668b6f01d04ec86fe3adbb1d10cf10a",
      x"715665e55e747c48a78af33d2b59b4a311453eb4fa74e321520740bea88f7c08",
      x"f31557d55bbb93a1eeef7b284fa7d1ceb948bebb2b2d9ef1eff86c74f0bd8453",
      x"d68e4541450aef683f690a905dbdf7c43b4d9b99110e151c056c516a7b19d05d",
      x"aba70064b8d098bb079ed051d200d1c84d5192392d8a152928d8988726f486b8",
      x"f8e117ef071e09bc7d933bad63de7e9d1d98bb206581945ba5c0ce00251678c0",
      x"5cb25de4ff3db416c1ccbee473927e84102986c21d3cae89cf5c92dd4355c6b5",
      x"a8b32e6043534d46e77225d29d8fca0166f6c2d5aff2a5b263add769784ef684",
      x"0848924da4b98e18c8439214dbee6606f2f973d248b777a3f26ccb96ef54e897",
      x"78009df5e01f02cf33d75301440333cb0ada901600b4e1c14dc34a0f324146ef",
      x"d697a1930b589a9757c425fef5969ac12b5b298631aff303cc8f477fef4d6b72",
      x"323507a5090fad08904e1bff3996c1b51ff162fef82aa5c1bbf7f3baa8661bba",
      x"b5f41fd67398bb4d6c7a75c73d8022dd55b52ff795b634407a9ea6ab6789e545",
      x"4c223d6e7d98fb90d6a6a5c273bc12d2966c0ce1e63948ea0aa680692126793f",
      x"a4335118bcf3d77784ad8167d2af28ff30130f180194d73d4f94cc1b9ca31aa0",
      x"03ecd484990f432ed325e9076d7585ee09a54535ea87dbc474fd0180affb217d",
      x"0b6f1f7fdb2437cf7626b345e71ba651a2c19e6746be15e936375b7cbea7aa4a",
      x"7c8fa46dff2d706412145a19266003a673fcbcc06d4ba58f9597bf9ede6bb02d",
      x"105ef91fe75bec193056780cddb8404198f3622048c974f54cd06f987fc06f9b",
      x"2c80a4abf899accfb8edcb8e6b98d5a3b1713fc3b63f1f249b4e1e9aa87301fe",
      x"8f13bf1f6bbf9a54c835740866683331a1b9397ee45648c808191b7941e2be69",
      x"49f3a60cadb226378270d98e455f668eaefb7178675f4522216f838beda2c5f9",
      x"3a03f8fd21f16e96cef27713f33a81aa23fcc44f471e13962e0e35ceca8f77cf",
      x"9dcacf1e54f55ca40203ec3f72fb4e8aa458cba817aeb458ae1eb0b599b66683",
      x"d911e505acdf8bc57ed7099892e3d856ccdaa99cfed7a9e5adb58209ec47a153",
      x"072be3b374e0ba419b833b66a273946ce3a6c9a3d9a9fdd5b266ebd14a980a4c",
      x"bf503fdb806f05585c69587b6c003d7de6649b312d36a477473f4a6eb3cf0ff7",
      x"751f00c67bb3a211dcea930db661fdd37c6601aadd1f50763d46a17859ee739c",
      x"f92d401eb3b77d0a14e9017a5c71633111077d811e47ff5f5ad466d4cf1df682",
      x"f417e5a2cfcc16bfd1bee4a16a8036c12cb0ac98cb841b6fd76e3f90da99c669",
      x"d2c186ae2f5a05eeb0b852d4e40d07ce746224dc074ca2b19e7421c5d3275999",
      x"661f9564d75898e8ccb1da3dff4f700b900afa22faf6d475e0bffa23eb3cf05f",
      x"6db96e956d8e0111b358c2200701dff9d7a7796b182fd54594371c6fd906e128",
      x"2971d08e3a337bc1fea5afdbb0ab37eae97a702b03b2f77f85f16424d8c0d476",
      x"f595564e80a434bf51b2db3836bef479eed7f53fe49213a93e4c274261510f65",
      x"dfc351733e23f82ca622c1ca5ee5ad24d7d86a5079d483ce415010cc22dec6d6",
      x"23b6f2256ba2b0a1ac4e35a0c10935dc9e664d14d1626e57767774f10210c5a9",
      x"e6a947f09584910b9b285b515ec5ef7fc0d5d41ed9332c251e6ff203631fc56b",
      x"471e9b0ed1b7a3ec566cc18ea7b5da261def77dfbcff4f5b46376277e77abad2",
      x"ba56d4e97b4c6a098397346f11ee547d22a3011e08b16b8e0bd9494c88d71379",
      x"07edd5426abbbe9d2a0b3988a5a7f95282201b367e715e6405758352dca9e99c",
      x"6776a1ef43e8e3b0a96467cdd2621d136c4c62dd7f91838afafd5212626d8634",
      x"530e9c8bfdf5a5049f6f58841de1f5217de1da44eb5c0051d96f4763586deaf5",
      x"e73d210a76eebab72b36dcfa8735e1f9759293d03e1fbe5e096b19f8d9d0d921",
      x"c1b6c2748f3ad8d0ae5206063ef0b95d834b81322775eedcaecfc932654468f2",
      x"eee387617721fc15f1c2b21ac7a0575c217987b564f980b3567d11a1a5ef2a73",
      x"ab06937ab81937a82c031514ccd6a507b021b33b210ca49ed9cd8b343bb77392",
      x"ac4e55feb297a0074a93099ffa811c8d885ca421c3bdc48b96f2eb165cc846af",
      x"c67921f8ebc2181c19f8eb66a8517ef39e8d93027888b22bef522a14775bb63b",
      x"654395cca07b96f4de5787d9abf33bc7eb2fe9327c18b71646793db0247b59e4",
      x"cc2211ef199378e2e8ef0a69b691609fdc7b7733cfc2cd75f95c620417670541",
      x"b72090538d6bd57ec184e0dda01886ce61daa4120a058dc6dbb9695a6df6f652",
      x"5498f45186440b028143ba5ac1289bb4ad408d7b8cdfd39d64bec07d38afbad5",
      x"951059a45861daefa5500a78be6724125ed4a13d571d57939b4c41c579d0f810",
      x"7e3aafbfdda1b08285c58486183df022bacd1f4e576a36c5d0c4d640f4b3e48e",
      x"391677a5752dd4f18a817c48415cbf0765f9dc1808a2d12781cd74f763d8ff1a",
      x"e6a3478cead0d4182aedd0248bb35e5541fd6fb68cd280eb063b1aadf960b390",
      x"a027e3fa1b16c4519abca262e64445f96fe1eed078157fb174e7c66edcae7db2",
      x"3e3269726b88c2bd387fe3635e8544e95cd726a1c175c1a69afcbe7a524decd4",
      x"eb4ceb8e1caa0ba56436a86ceb807d572a9774a6bbb04c1d15de6ec2afd96eca",
      x"a15277350f9920b789f1c9b0c848257a1dfc6bc39fa0a5e21ec294c53f09f688",
      x"ea3fefdab0109245b4b3c33fe5e2a1ca1fee4e2cd987482ed89bfaf8becdcdfc",
      x"f8e3da289039edd51423debc69158fd2ebec130f46426691bccbc2ff703469a9",
      x"49e9ea444b6184db1d3726d3907709183be813d6abeed9984abf67acc5137c9a",
      x"d83c3668c595938d1c695125bd15c8a0d80493906617fee06e34648a7430cfeb",
      x"cdbc41a8176de619de710d81e5c93e45a3254b6f249f408279974f6291aa7e06",
      x"cd4f62bb36963f2743c1ea2874c7dbb9831bc2d6ef14a383a68c0061b56e69f7",
      x"30157c38529325d731ef8f55bbe75e061b2c0287a16a046b1a666b1684f599cf",
      x"ef10517bb619c02422fb67e9947cc7e9d6d5d08a6202b29e3274daa073b08c0c",
      x"180b7a61874644c514ba64858a5701fe23de9fe3499d286b13a48c574eb6c8b8",
      x"808c3bbffc31006d531cb1a4f9736c8d03f6de969109a13e1379190e540b8523",
      x"5eb5f2f3e5f2de0243ca46ea056549f376cdfb7fbd66c2376e75579f071e3af7",
      x"28dce7042744073078ee50dd013aff511ff1a7b5c7314263892871b0afb2d22b",
      x"ad76fa30be163661b2d14943c1119eafa2c563d02962d838cc71a4db2b4e9a97",
      x"dec6ecb6b9273a0ede5d30d59ff5f229dc180fb187a342d8536ad05fbf6dbf8e",
      x"bb482685a31c1d9891d8b292fe7fe7b62017f1d8123d1923aaf4ec6f34ac96c6",
      x"a75d8a9a3188ee8698c31b227355f0c3fc3888dcaac08de8baab22510ba77190",
      x"bfd4ba0b2808965dfb3a7e9423fd52d1c9a7c98b656cfbc75966af9eda7cfcaa",
      x"9385c026dade442723f2a0ea0e8ede38aa0f5ecc7a7aa504b003572fdddd00d6",
      x"6f550b18a4ff33c9028aa629a9f0d24572712c6617d932aab3f4c9f073170069",
      x"3e3a7089c78c9ec2ef278ada7a116332c0929f5538b87fcacd7dc7a2282fa33b",
      x"096c6c05e5349d09900e4b9907036fd993a01925b3fc5c52becb4567ea0080ef",
      x"b06547e358d37f57a835b77f8e93a9017824f25690a1b823f14f23cee3713ba3",
      x"6cf8fccd73237b60cd6234e9e406ff8567c094bf0e8053410eea111351620650",
      x"c0ba772452007ca49b88a4c0e1fc54fe45872bc1e62b95aa45b88c7eca285c1c",
      x"7e8397b953a248f5fe1462f751d1f4af27ce523510e93df39318d979e40c2d59",
      x"ea3fbc7cf38a40cbba1b2c4a3913fc1dc024d4a4557072940ed7b0620e73cd79",
      x"f66ecd9fe5a8dc898340263a32403680572fda4cbbc266b55271b727f87eaa94",
      x"7473a1a378676adedecf7e7a2c98db49ecfe2627bd2d3d6dac1b40c175e14390",
      x"c46d59d847a2ebe346c951ed3f14e05c2cbafa072411e3f20e503f244639fb0a",
      x"7c48377d4a82ee0807a7f1cfbd9243185bd19485b1942c093df7f67d1667f45e",
      x"ce4c624aede20cc15b3de99b075c5e4c05889d61d75297cba530ad9a80682e99",
      x"d8753cef662a756390c26ae4da433257bb2f4ac44cac31626b8c394ee28ab5bc",
      x"018788c9c72609b5f153b9a320067b7731335e5fd0fc3d961743df7889cea111",
      x"2b721e8170f90a9b31a22b9af0d10e823b6d842f541013f8741ee9228879bbeb",
      x"2e1ee45284d8f1b07677b1833c899bca72ac7475f7b10f3109752061b16a41a7",
      x"f0ec1f4db778c69ca967d4a6d45edde5e0698a9bb2184d0bcc4d752a2bbb7742",
      x"e68db5259fd075088dc96e166e85ab0e1c38415b5746d8bc4e9faeedf106afc1",
      x"cb389f8b89b4ea86d2875821f3979d677e79c0484a6a8113eed1101718cca95b",
      x"cc7b35c99c4df367cd6b8cde022ab4282a6847ed81e6dd2bcfac7a54a98d1936",
      x"1833b5d49546846fffa3fd719564798997ed347397003e66284fb67a63e0eaf6",
      x"c4d594cf7a75ee9919c94abefd436670f15ebb34c32f7e121aca27a8fe1b5bcd",
      x"0eef8db2150150899085fcbe3c1a23d48e8325131965ecb3629bdfcaa892e67f",
      x"74a4e1cc8e02585c672bf6dbad110a7a633b6f33dc69870724109c085f378196",
      x"644cc4e94385ada2331ada7e2a7d0329f31e8726dd9a187ca7f0d07824ff48f1",
      x"1fb2da8647dedd536a9fc857db6513285817e0b06b24432bede94ffd816ef017",
      x"58d5d8fb17ef775b8682bc1ef68bb2d6bc6959af2fed2343188804a8a0b4b087",
      x"79e8475a9459c25d8481e79075317c408f20571003702692046081cc81859de7",
      x"6bb6a61a541cbc3cf4267327df59daf9fab5f41c6c79366671520d892c38b8ee",
      x"4fd9a274361428350b9c824a431dff7ea18673b24de1774891cbd88075f86208",
      x"4d1663363dde83d834d1f0d69b9499743d97e85a40592721b9c322f7a8c42020",
      x"7d411bef46863c4aaa1a828375e72bd7040a860dde45973af5059bb0772c16ad",
      x"7c74a951b7b82d3a77fe5bb15b1c7efc9e0c329200d9ca1d6d5392b472545cb2",
      x"68e5dfe43bb77e66bd3c6fdc8732c49172fd2f35b3350d4b2657ff91d182bf87",
      x"96c850e217e71cdff17aa0e3e2139f9547ede31cef91d2b10b53058bcb8fa2cc",
      x"374a0bfa87b4bb599919c85d1ba9ca028ec022cba6686e03fc09cf4992fcf3dd",
      x"be1d1ebd1828f4542c8a6ca6b59b0bbcb4ab78612c42a5dfb4b3ddb0273fde71",
      x"dd9c42a1f6a4c53bd55adcab9ac7df3c8dfb9030a8fac8dc5abe93289a84a429",
      x"be13243f37c528624a3abc97a0f0c9f4ffad3ec6ecd142df8167d42fd55088eb",
      x"350548485683a23cef094604b03612bc03be094c8a707b75950a951592b96817",
      x"b4f9ecf5d15f3ff5923aecc610969e5a3a4f1f6834e8de68e360a5344ff4a363",
      x"b715fe50f03cdb43242ef506c7d98fe3a561e21e0c250d4d95a9460f77267442",
      x"6dd9e9499ccd5b52f1c8bc8657a76bb4edf45b37d5be49be6be77e6e65267f61",
      x"fada5bccf70ce9319e9539a7a720ed52631da34ca6e3cea634f3c15275448c43",
      x"99143190e5aa62d9f8b4ca591843a5fb95cee9522b915aad50a4762c89d86480",
      x"59e417f2f61cb0273f032496d7b03817e241da681fc1135cd23fe95be60ff213",
      x"350f71f5bb7795bcd1ef937bc3c3d74250bac5ba361142abd06f5bbaa42d5b9c",
      x"03dac6c9f4dc0710fe79d22ef4e28ece8016c92323e1a17e147ccb359e7897d6",
      x"6f283d5a20b41ffbe13932bf15fd8b804900b1b3af674a0cefcd817b04f8a2ee",
      x"012a192e7bb65f733a4e982350c8e1c3af5ee9f1e1f9e8c50cd379f8f44b0571",
      x"e87b8c1a75d2182ef0dbddc5c944413c06b927cce18b390c0d15ffd2e61ce662",
      x"44e0baf264362a85f2ac6c24aafe41a66d3795535163516510ac169760c2bd1d",
      x"0cbd236864ffa954b8de523b4c3169628fd447f52bad2e0814e857560f4c0752",
      x"2f92c429ccf4756abb5f928af9a61a6c04d4876b57f2c7abdeba93cf3b7d5418",
      x"b7a664495d73896cee0335eb5ae854da32c6ea11faf7f0b074dbf2804445288e",
      x"c3e643be99ec8d951f2e1e1d1619301b96d0b7f4fe32e46efc3be591e8e9618f",
      x"09462b9fdb948169022601f7ab5c43c98a61f20da4724831470f1ff3a6ee6b16",
      x"9e67c2031724dd36f099bc15621254e91000d9ad0e9403550287a0eebb0e6c99",
      x"ac8c8807decfdc760a65395379eb5cda210bef2f202ae5c9dca88f6ed31e2db3",
      x"6610d61fd0c6cb37a2b1785e6df6128f03788f59d1bda6ff7775d7287b35f7e6",
      x"e769e5e18eaef81d152cd2839a6737c7b22b255792e34a81366f6cf0bbd02dde",
      x"316dd9e38c13e4986d0e1dd7c1afaeb258b42b55469b1f14f13914eef2e677ae",
      x"43850fcec7968ad9ff0cf47ba3320c139d988725354db3d9eb39d2a4c1c6111e",
      x"258e0baec9a294adac009eb1e8e3152dc0944f63a08b231a7f5a0d54547700dc",
      x"20b6431269e272bfb395e75de94c85a786ce7186615214583f0f803c38442a16",
      x"364bf2a50b4ea26d105f3c4d898f5dfede3284b3550b19e175176b13207c29e9",
      x"b6ddacaa2ce37638266c9655dc98b4e771847937f3259a34362426181db528df",
      x"452f30bc11fb73ac2fcd42b3c28dc1bb55bea08dca0dbd8a3ee74651aec4cf16",
      x"265ed2781928b2221001938fe0c95621db7368ef3755f0940015675a826b090d",
      x"eac39c71df0857b548f94762a038cb16e47b0d1a15d844974c255bf28a00f611",
      x"7a9d290c63f12de4e643a6593c826550ef9ba9e6d20cd24b26a722d1f3861315",
      x"6eb4199fff82bb262a96888a3907a387c722802987dec040ee75ec0e971ee9af",
      x"252f282769109bafb4790a8f24bfe151ab72ad996b0aea168e4a4e7f092fe134",
      x"807bbdf6ba18a3c4919892cef575a8c4cb5be5bb62f687163206f457e8e4b6aa",
      x"ff94535f4fc3282f867c63c3cacb8e3f8d915476c24f76a189e3c7198c24bcac",
      x"84dbbcb181fa0809fb74e4c2e40fccc9deb5484a56b877cb764b82e135cc7e0d",
      x"9b61010498c4ee73500865a092ae1f748af89dde74b8704741d6d9af72e44a6d",
      x"1e667172bff6297ea391a2f0f115c4b53c6d69b4a907e1d3940acea9b7645d51",
      x"c3cc7d928c84c454678465edaa91bfaec23122f6ba88fba69c7e5634aa2cc00f",
      x"44b452c755c20200b66fb7e8fb307c1696280600566aa3f598e37485691e4e7d",
      x"953c329f94959f571160461d39ad50796753366a9b87883204a80fbeab26488d",
      x"15581d7fae3346a371fa662163fc957cdbe7f370de7a0dbcec71badb0a42e13d",
      x"64a913f89330442f5a92b26a29cad8207adb8d87a0daf83dc4156f3047484618",
      x"e006e9cb9ac6912568fe3241172ec83e7d6c34e65dfd248950958f10efc7177b",
      x"6f5d4d651a4ca70f308329c8c62e1e48338e70af226160ee00709003bddf9df9",
      x"39ced9bf2a4104726d5a033b50db6ff345b80a74bf75d60131d6872c1e2ab5a9",
      x"7adb032b53f397336a1fb8a325fe2eb81f87516f05a4cbc1b49402c814143f49",
      x"b11807a8806c99f35d47dea58094ee78e242a474be2d2cfd686cfeb1a3bcedeb",
      x"3d51cc88c99f6c5ea10c865109f0b0c2b6646a5c5441f3f432edb9ff8d446a6a",
      x"7f1e623a5ea543ca68db7ea91920470bd900d57c7998c8bd9fcdd9baf8ff775e",
      x"e7a79105518dccbdae32d4558d6c7fc2b780e0202120204af87af38e6994c271",
      x"74d8b27a11753a93a0275a2d232b250fb635bea2a88c45f13523b026cd51b4d3",
      x"703edc6623563b4525e94f01d4b3bc128b706ad1586ca9a1da77f28ebf8e7774",
      x"ed41bff2717d64e41474c362d6b8e9726e6c2a006ba46aed2c9542c19bced857",
      x"f9a7837445e6ca50b3487ac4d71290d754258dd7e33bd798188c82d96d8c1676",
      x"8b0648ef4c398584ad02c2ef6c02cf36f21ec66d3a4dedb7413a6b9070b69eea",
      x"e144d543fb07230fd84cd1a219a6cf4cbb0eef919e2bb018e657f5f864a4f4a5",
      x"d08e0b7a1449dbde12ddf9c27d69ebd6ffcf00b325d854194602b5fdbeaed573",
      x"b205aeff1ee15702a2ff55c4a50b022ab92b7bacdfa37683b3b52c8fca357f74",
      x"50b8893da17575ca9c61c5fb1abd4646595da345623993b80750adb0556b3d15",
      x"b59df68bc8b65b310f805432ba376d8d8f901df537b87b6570ccf5ee70f8ad60",
      x"a9ee002bc20e7518762535b7fd727b089deb827c3930d46e3eb6ccca58111f64",
      x"374ed5c584ed4069e614bdff511ed0ab1a027ed2e422dd162852ac4fac026701",
      x"6397dcb1c9795e2a4f49f5b0093820a0525b71147beb37d4fc35c0d71c5a30d7",
      x"71253623f39896c94f05ed9f9285e9651a7e2f95a77bad1c14b345b49a102d9c",
      x"8d6416e2d564224e337babbdb79693a106270c28a3dd04ccb7283e6da59ee0a2",
      x"0946a566f0b4f5454dc52793dd9cbbcd2cedabe2316d68af11f0bc3561c0d751",
      x"3dade91ac2021058f23bae383de865ede4ed7a2d51b62acaad08f959f5da0166",
      x"35cea6ff43fa3089deb95a4db6328c19ad3ab1162af1675dab5f12e04533f224",
      x"6836062e1d51cf071861eff0c677537a8d8100d7d98a12b2b391221ead85682a",
      x"fe45998fd062cc8baa3830391d6d347a0be1d6d5e05709686719e43a4c725c9d",
      x"b4b17dfe85bdb014faa301527c2601e36eeb52b5f13eae2f3fae2449466620d2",
      x"a1ec7b3e3ee8f9521475ec8d18a13e42c776ad12b1b43a00b764654c3ad31343",
      x"e4016d3c2691a510053ebae5919f0f6ec056701c80a2f1a8f7ddebb7f6fab57c"
    ),
    (
      x"ee7d19fbb24a518a0e70cf6f77e0d39b0a9cd260fac582f0f55ff8e8dc3eb9e5",
      x"77a611672f1c455131f1947ff54d9c65b89f0dff66cb302e085db10516d0a31f",
      x"c7376abec801e5b87ec4d025021bbe4ee9d2eee45995dc27466443463e8a4124",
      x"07c83e035d728742e57cd9917f7aa015406978738540deb7dd78edcd3ebf29dc",
      x"e30a63a0325a7b1c186465a534febeab29274c951afc98a73f8b4700fba62d35",
      x"48588cc82f5da7ace328485f273d6d2fcc580914a9f07ea984bba8e7137c940a",
      x"158bdc5a5c7d8bae09928855aaccef5ace2d3dc15770dc2db90d1c0675b3c3f7",
      x"34c550d4b24b05dde9e5327cb982138fe709a785c529491531e3c4be4c8ca327",
      x"bec2ef38325657bc28bf3daa4cdc2d0bfda15d2df8aee561bbf4e8fd34a9fc47",
      x"fd9ccf311b7e98398a8560eb430a626120de82501a475949325a8b636aff8ad3",
      x"fb60d141c65822a66af679b7ffa40737f2fcc3d63d6544b8684a5e2ec0ab739c",
      x"da6c58585a20abefce0d0ad0c6464eb71dbe0dcb87d0d5d2cd1daac8848337ae",
      x"81654edf9f56748a8f51e7ababfdb1add3b453307db5176599f1da430ad32afc",
      x"b39e6898788d6deca31015c891144b311df695a9c40ee3563043e2d8fe96d8d1",
      x"8fca7364f74a1dc72c56ddb891f22dc09a5dfff5e9583affbb19a24786505d73",
      x"0bc0f75e7aa00f4eb0b8f8b1f210baa5376047aada1fe910b097b64357911560",
      x"f8389ae1f5be20ebba867dabe33712f1765ce1adf79311c78859a1762b0fafbb",
      x"2303f7c2e190e506a761fca58fadab96731e9194516922ccaac4e2018568b9cc",
      x"d81994a067a5aba20f1980fb9de90ab9caf0eba7fc93e8c92a0bff713f61cd6b",
      x"4839c792b783bfb9d47d42e809a70cbd96aad5713b11e2fd962fcf638570fdad",
      x"f901a14d39c06f8106e455001d1c6dbd0bfa91c151ca372b2d425c3a40f21e41",
      x"6bb7a2985955937a5510ae25f79d391568a4baa58a78a43e306e880f75fec5e2",
      x"166c3bca8068087d865b8557e6462993e7cbfb6f1a4aa5c87d0d0d62bdbbd6e8",
      x"1f6f2c0570058691b67f301641d599f7a78d93c7baf959762319e6c8691287b3",
      x"08f5bd17d6ed179040dd7f7e5648ebadbd99b6e16e915cbbfb32d05a9d297b61",
      x"eff4f8577e1b4ef853aa803cb6fd8d087ca51526a5bf60484ce2ab2f4c66ecee",
      x"b12ed5e6ff2a6eddf07c6a13ac20e6c4af739263acdd3ce6c8bb03e7c9c16f7a",
      x"18d0aeb8a89fc838f487605caf92425e0a1cb902dc301254604252d929379e81",
      x"927d9254760751e0d2bb779e196ed11803bd03942c710e94fff10c40b5767e7d",
      x"14c92193361f4d59608b614ac15a88f9d03f20ff880da6bf8220e744fc34ad01",
      x"a2f765f06edc5fc4f5525b5c1eeffded95da681517c8bf924a8806fe1c28343c",
      x"6f301d072b5168326f5f30bfacf5009d82ac0c1a34f9fdb8308dd29fda1cdb14",
      x"bb31a300520d52e5438fa7dbb4b6205109c783958ca932daeb7f0527efb30cb1",
      x"4802a17467434ed4a3391d89701c72ac543c2be0af6bd924debc855c9cfedd68",
      x"379c4ac0005be2b843d4ed7db86c8c93790ed688bf13c19534883d75ad8c4e91",
      x"ae4e23998d22bcdbd9fc839fc04ed7fddb377f94a686b9b9711ab8fa0449ab5b",
      x"14c8e2a9e2c9d3c1d8cccce57f9ae6bab667ec2b5e9e0e589342e7ae58ceb596",
      x"510f12c0e74945b2d0820f8a996a983ece12be443cca068f7cc5c211f57f5f68",
      x"e7e52aa4ce368c9e8e8e6d9a5a9b678d3bc670a93d85a75959313831b36af5d1",
      x"343a8047bb2c6ab3cf4032b255f21dedda4ed986f0f35e23a32de68fe566da7a",
      x"08ece5858b25904411804a25a790f3e9ccfebde15054577f83d1ffef5992222d",
      x"abe50ccc7006291c7eb23edede176408cf44383dcc0c00a08c9deda5a510412b",
      x"e1a06390e689b7f5579bf4d75ca000f74aa44b3ae506e966323fc979d6d65966",
      x"c3de89bc35633925d5633cd6233f41696a1630303d42b0e64186f4cb6e2d3070",
      x"054aeb0bc147c7a096c3acef03fbc62add37a66f6faab89b0fe4db0f541887cd",
      x"f467de4f30e726d6652e5f39c75a235e4cd6cb4c4044f7353f64b4c13a0333f0",
      x"6cd942766937c0619c617f1705741d21758899cbac537be55e921b1bd03f6517",
      x"202209120b9c4293817d2ff9b712f63570826a2680ceb5bff5761400237a1a6b",
      x"64b1853d180ffd015b9b8375916b195956435abb6cfe392631d6aa763b029a37",
      x"10c12ea54673ed626084c52669641101f81607446c019027be894d62a52dba5f",
      x"26cee079e7d0ee74f9032b52d1710c9f999463bb2913fa33ed096d1ca3d1d071",
      x"6cc09ce7402178d14f52bf39c148c1497be6a791d0b077cf5ca0c3f45fd47e59",
      x"ef7ed4fa666625ceedf396ff2a751d298af38f819c3ba8ab81dbfd16bad9358b",
      x"6ce414917e629467f81e5bee8fbabd1443a8655b5a5c5d381b573f9531fbfa4c",
      x"ca762340155911ece090568f62e37c9ff1555ef95a0a2f42dee8781d0ea9c871",
      x"7b6333436680a61c431ec8880d5f2beb470e1de61a4f8b7ee6e3a650db07d792",
      x"53e41d680266525076073e462d5a962e5f4cad05d84fd87b02fc12a2966b63eb",
      x"5752c69fb3b6df3119206c7e874d6e32799e76ce9993c27f26fe997dab6146e9",
      x"68b2c4fb257149bf22f5416432b1d2c9bef76ae0747f7751f628699ddf501506",
      x"c272929b795d9bff65434dad11c1c48f72defd42317d98dd6324958babc84c53",
      x"62c575aebc732b706f02e8d69e55512c3f0720d25ee9c1ca7a4ae7f4fada1a8f",
      x"47361f98eff58c1e37a9d33b6dc514bfdd3ba69ad50b1b0a817fea7f3907bb41",
      x"e22c614f61ccc76d044aadab24600f14961fef2af68ca78b543f3d8420b89435",
      x"046c16b80c5378e9956242c9f69cf3fb3a60fd63e19ba4f6efb4f602f9997fbc",
      x"55af7a9b040bf91b0bc9be18949270264694b93278f87d9c86bdbffd907e75d4",
      x"3677be78d01e0a83233bea662f0ce2c4af86f97c6a13eabd56d1d2b177edc8e3",
      x"6fb79a8baf06d08f185bcb982c4db5fe82abb236b438e86fc6d59fed589c5d15",
      x"7578cfac001bae37e5030ce623c2289483f6a8b5f655a0f6de77a11a18755d3b",
      x"fb97a9884014a7ec440bb2713589d3210343ab4742597237aa9cb8ced8d1a1eb",
      x"84f3b6af5c284e997b435a5378070bba21d89c41eddde7278068f84b04e0dc5f",
      x"f31b8be80873215390ddf41a1aaa9751c2fd224be66fdc48e929d6a093db3bd2",
      x"d8e9eff66d8de27652acf92cd4066703a6432eeb277fae45db691e213ee620a4",
      x"a0c040b92dabc8439347dd995b1c20ba3b8dc82d723e4a70dd0ae7827bc44ac1",
      x"d7bf6fb0959c1ce6b87d07b505afdca56ab6bd794a0ba97a6da32f3c1edd2cd8",
      x"d94ba73b8c767799361f9ea2e1dbc2deb3d49203fb0698b75e266ec7a284ea33",
      x"b50f80134ed272e5d660d9c09b2da151dc026c7c6cf1ae0ba545ee2acec2f2fc",
      x"67355c069f6936e687462bbb052bc0e2b131d0b217216aac29812b58e00534ff",
      x"959ac4f04f123665ea89cbe7d12396af138af394a096ead337bf4897df788bf8",
      x"44fb1ccda557a40b9329878a03d4fbb6ca55809db334dc137fab7bddf7e130bf",
      x"63060fa30f1feeb312a831db5e0e67adaf80b2c9d781f8e542681284a0ede1c7",
      x"3b1d24ac7cd987fdb6de013f888d916bf124864cabba145c62c992c2ce1db012",
      x"9f4d1d072a3f601c7abda0b0d3c305e9f4119d0f1b1669618602fdb43a3271f2",
      x"97ec59430bda7a9e160b3b50f24141d443f6d34d5ebef4952ed123a6b17f913c",
      x"0fb6c86fb260c3a35d9bd6aac0ec84cc65df45b350e20c73db34a29e8642a6eb",
      x"e9decad1c3b92e1049d86abe29a9fdba31b3399ed97a8aa8f3bed614eeea6749",
      x"f1ab5f5403a45742ec306cdf3849defc455656e75baff02b6d84dbc70e89281a",
      x"5318e296faa2f2a92b4c28db59572b7bb6fe0aae9b6b2b77bd842ae5144aab6c",
      x"1bcfafa6face55a3230cefc1df4a2e5be27180719adf97ffcfee87a5e8daea1d",
      x"98ffb60613ca9f7fde37352feedd8559555a3f19456a26a15121e871e4a7044b",
      x"260dc0de44110a03d521a5a9f7bbb1af57295d2358db4e6fc9ccdf40b190807d",
      x"341145f01836b27f09308a155e3c44c5117c4ae96a154972c7a40b2d226517c6",
      x"4c62564095d7fed7bcce46691d7b98717ddf201956df5f7cbb69990c3f976d88",
      x"89efc9d1d98bf2b1f68b2e42a60e4958de974b727c7b4012609f4ae8a083c985",
      x"77af6ed80f436e5b48e05ab7da0afd3b727ffa44a925c1d8b868e02225085851",
      x"1adc7baec21aefd4a64a057c3bc6124c42da21a2a9ce548d1f03305276444d6c",
      x"b65807461855f1cea7413262bf49bb771c9f6b6dbdb9bd6837193728fdd64c7d",
      x"dfb1ac89fc7233f6971a278ffde0b8fc9f33d5efc8b87eb3afd1f660c9be1092",
      x"259c5529e09b332734311e5ef192678120cf11c3840abc00fc39235b99cc0953",
      x"4165c40ce2659eb05b6205ac88499d972db9c6b32434c557a66c0a25787d89aa",
      x"e4894dbf590a353d9041f59877b77c552b4baa458da7fab73bce1e8f40cb8481",
      x"ab0239548aa737f5c5fe8481d02d5025e444d54e37347ed220f28ed9a6070f0c",
      x"36c387f94f109c512d43855ce4dd67c31f036f9fa8d21ccf29297c3c962b33a8",
      x"1b569b617246f4754c1378630c662bf4227fb9a292004663df1d8d1e436efc59",
      x"e14f1392b0d8670d31d966fb85b7ac27db095c1d037fde83b137056c6c94f3b8",
      x"a708b0d3ddb76bd78039d9f84aa01f989b5c24a71fe377eb114eda234add7c7d",
      x"5ea995d137a1d0c619d063ee44ed96165623b97eed963989d65431da904df909",
      x"566a8c7d6738493ccf046d42a3af67249e22eaa68b6dba985cfb247ad1160765",
      x"bc43cfc6a206caae9995ce3647877279f8a340def77a8c8065ea4d1c28f894cb",
      x"af9f49a2d8cc4691dd911f7e720f7763b2fc5cff7827a8dcef557ff2ba2a0b8b",
      x"97182407d47e6329bc52a8472b90f01abc800ba449f75755a5599a60edbd9b8f",
      x"606cf461c921e45899905829ca9c3b6ea7e7f3a77b2d50693ac67bddf72f74ca",
      x"83f1ccf3a13131cd9bd511050e0b09ecc118fad52275c60d1bde35f97beccb11",
      x"05c022cf518cb3ca08cf15cdc9e1180da8e150d1f15991c23d7d2dfc701f0e9b",
      x"137a9e2bf5b181f13ecbee4ef7927cef8ea24b25b2ee54bd1594860625074044",
      x"6941d17385918082a6de95dac31d43f41f49257832076505b4d4d85454211975",
      x"e62094a847d093f0c050e4a62ae2659fa47fa03b3ffe32f4e769b3e0237f9817",
      x"1cb5f868c37c1a2d8b3632f909a59eafa030f0dd11781c8d343f33c5b000b0b5",
      x"55554a2a07f2eb6cd232e14f452568f00e2edd483a27ab0e25e4b79a6152f4c0",
      x"33f5f576bf698e9d771821a1ee6e8b4e4b6007c9b6124ca80e9cfd74a5104248",
      x"1e477e4085fadaee458163c7f96338f6db64f3630503cec4cb218ff9485a9237",
      x"8efa66672e11086e17a8b55b36dada493c5c58357fb5b1cf964f39c16c25dc9e",
      x"4910ccad06f63caffc634f413172a859a90d4f05298a83ec371e3e128fec1230",
      x"9be79874841372eedf433b69df4531bcd69b9319853f1f634a71edc367b64de8",
      x"6976babe77d778ee012e5d948c0fe25110ff634d911dac98803c13c73b534d97",
      x"c2a0d8018b170f0c52dcd3548062d6500d9aa5cea68788c557822c7c656f7066",
      x"cf5b9aa0a8e4de1379751c5a24593d5b2c49c47179033a40470b3d10c38c7802",
      x"0e1da77f6cccb9cbdb7c8e1404f08dd1ab1602a2203229ed3c0cb454618be92a",
      x"71e14ebdf0e0b5ff424a7c81b222afa86a27ac0f7e738ede2ae405a59981e81b",
      x"612784dbfc8cfa78ddc024b2baa244c3eb475a2a3e19288132d5c85621d8f7ef",
      x"4791afa3b66089eaae37f8458e68701ddfb2e6d2b14eb4689d26bdc2d66b2b0a",
      x"5c5fc1611df3c4e34158bb21377cc09b2518cf741b34d781c062b1c4f1b1a824",
      x"4018a6c30de8cb4dcf512c6016718f581f2df14594fbc3807d9924e46d2b2319",
      x"c8f5157e7fe120efb92f9f7c6b04d56f5128d0e90db9b5ab0da40ab8e4595ae5",
      x"0aba9e8f96b6f246953c22c37a5c97b8cc236da7b7d959a5480e2597b27ebc19",
      x"f372686896a155933213450fbaab95d8fbadffa9185747ef1cce255b410c88ce",
      x"af73de9f96fbb6540528cc9145af90ca786fd073718f6c900d83cdb0020d18b0",
      x"ebb9748197e3a6847e412817179631cf4e8d0b6625fbb9cd2aa4bdeab507b2ee",
      x"e0146ec16c224349ddc60f90f74a51aba60fce18ea8b2c67e5062be28ca19bc5",
      x"ed79020a2f0c8203e4d4283b66ee863b7ab9c0ed6ae39ccd0367852690d261fb",
      x"30fe063160341cd2858a2e1283a160e140bd82153e2d48a087e7d34ed5fc0b2d",
      x"d20396c738b4b6a0d6a786d18ffe59eddef524f55b56772939736c21fe8ec20f",
      x"4ae68fe5cab9317df1afaca03d0e58e2f4ddc1e5ed763411ee6dbaf1fa3263b6",
      x"ad6fe864d90665b9772e39b629b1ccd638fc781a333bf626edf81babccf445de",
      x"77720df5fa48a46ab4af83e7024e3a1c6a9fca3946f722fd5b0c1198e3717538",
      x"ab3e74450502bc715a16de77eb6a87458aaa7fa80b856936f83eac2cdc5562bf",
      x"8679219cc803fdad5409beb6661065b1d0ce07f648b5833622d86e9d27c4c372",
      x"9846dcc2b1dd0f8978b71b4563de6079b7076589b219b3f7ce945cd7c57167b4",
      x"330d41e1e96681bc586f14bc8ea55ac625010c7132b502ca5d987f7174a820a2",
      x"53792c7dca136950736c277649983f5934f1f8647b551748d960ba86b64c2763",
      x"0ac09ed3c1fcb63dd6fc7eae6da512f2ca27c1881b32612270398841f6747807",
      x"ce5ba62ca530d873c68bcce2057d5355491fa3d8b683828c26f55474227709f7",
      x"ccdb7c02af82e080817987eda5d06f3801396f17c49dd29d32e6ff0205375ae9",
      x"523165fce83ac3cab5c6c14bdbde7003fa48d7a35cf58a99dcecf35c753f2729",
      x"ed1e46e003eaa2b20e746cc23d1bb7c2764f2709e963ddc550e47cd77e31e0a4",
      x"836e741890986e032ce7769edde6b8216fe635a1fae087878f2147373ec7744f",
      x"f9ad876606382df87bf172b27348402d7ee04ca42ce42c4d262f80f4032d749f",
      x"1804fd721dacc56783c8e4f5375629a3eb2277a2ccc5fabd829734304e4b966e",
      x"502cf2420e28d2f6aa50949bd3fd2c0b46817a71116919f89dc8fb5a88b8942e",
      x"e81211876be8e2c965397fbc19e3acece97e9a1ca7e874ff8b3269416a613350",
      x"bd6229869172b0808251065218103315aae8c927d07c1b15823f8aac1fdf1c5a",
      x"d3528d5eb59a8c6ddf55ec6d5a930ec843560300bb4f4b1463aff3dd14718807",
      x"7583d6b7c4e1ee735cbb426b9271865bb81e20076e5524523cf7801bc9db7a4e",
      x"cef7e5d38b9771c24c5f172729462b22c166a6f1b699be5bd1f3ebe373dc7fce",
      x"907c19dbf31edac5de08ba89f19595e8f8251a628a205009436ab4c918187730",
      x"135ccd29653a9dc8ad9c2d19826604ec1e9f86853182caa2667c634e3e900507",
      x"b3e0f0cff175cb4b19341b62dd2b7f829ecf5a35746cae70c3847de8aa7f7879",
      x"b62e76e3696bea5ea4ca2ca40a9137a7c87728a4c6f500347709da9a4ebb1ef0",
      x"16adb80e2c86a6cb74a5b1d76fded60637eee8b8849c431f18cef90a2d6020b2",
      x"3f4b4e7d5121efc99d113ee0d260ac8ce5014303fc0e6d986590bfb5bb9c3142",
      x"a5e072620159cf733630f7d98c89ba2939ac4d5b58fd1dadef8d3f5968b13678",
      x"564afdb0534167bd2dadd710f26675f0dcbabe99019111f1fd7dcc9ae0d29752",
      x"40d4f55500fdad00841729c3ebf356b26eabfbd436c33701f8bd91cf6a85a4b5",
      x"71df1166f90180938e8876b929188ef2b8abc2c1cb5b911e7ad540ac281fa055",
      x"b45ce06d5195a30f15e3ab0eaba1c555d7ac0c1828c552f2de7aa9a0e893d473",
      x"ed58d294cbd94c3a24a048975b6916518726722d7ce4565a01c8b5019af4f80f",
      x"3879901054d14e0ee8933fa919e62cca178589709906b16264bef7977dbf3ccf",
      x"e5177fae77cf092d6f8497f0bfd0dea6e561ab60fcefa061fd80044cbac25ac9",
      x"db9c5eac2ff2fafafe0a76d6a95afaaab84204e680d16731fb5bd668380fbc1c",
      x"eadc54fa6a6fa313e664e30f13c326b04b1436d3a6dac72458c283acbba44bcb",
      x"1260cfc5fce4ffa214b0efd40ac2ed8022b6e8c79783b1c214a4175a4e3dcc6e",
      x"0c5ebc4928411056a630b4954206888135be6a5a40b713418f9f75328e1f4805",
      x"2f29790911a026ef3f84e7fe141eb3d78f804b09e2afc419e47b5f46a18ff4b1",
      x"2c7b7bcdc203342648110d3ac3ba4d8d49971c687a6a55078cc5300d4b4c6a1c",
      x"be5d74cb880b15e7ca9fbc835b9d31a805e9a195b7df3386e15ecb30cdefb091",
      x"aa7ab15d10757990c1ad65bced534b71f2909f293465bab34a3fd70157897118",
      x"36d856a8df06be2eb760c70afe3823e4e4d3e35995759042a1a0aed8929ce067",
      x"1e2fd937bed5d5b8d01232eae86ccd17d70be6850ff463e8eb8de43d46b23396",
      x"9f46cd57251dc27f2291db755c1497e4f107dc922e33c0ff2443eee284f6a1a0",
      x"87a95dc3844db3d2ef1aa9293dbf88a5a5bf396adbf2834e85f137d0ea677ee7",
      x"c52d85d4bebec6f2abb4f91145153c68990aac0f82b9c25f78278192ecbea9aa",
      x"15ab4aa2855541f55eb124c84df9ea4128c20070466215e7edd39296c98ec15c",
      x"f2cf1e886c826557b4cad0e552e0c02d1b2702a9289b5af98193eefb0fab318f",
      x"df4f64cd4d6ad88a31481bdc560627c6a89a5a34194cbddb14c945a5de0ec911",
      x"6bc8397134aee0ae63f69cd38ca63786579fe2587e71996bf3fabd596878363f",
      x"ab825d94c362ede3975da4800c6936a8732bf0775e482ce738e671bce9885b92",
      x"1bce26f1ac736767af94a584636b5adabbf5c27d30dd22aa3410ed5a9f390fab",
      x"26296937e6ba48981ffeeebb9945b7a03d91d45e09c1b916254682b7274db4f1",
      x"8b752f46d0df00106891069b6d419079af2502d9cbd601974d48207401fd64db",
      x"5b878bb3e72dfe93ad275a2dbd45679f66cabeb55e8695bec2d398e0f6d5dab2",
      x"65104467cec25f35e3e26d322131bdae1bec2339062b0fb7863e2a42b853bf8a",
      x"cc817b3de41c6d3697114b95cfb0229098247baa5c46a0175d8a1b2d1121a5d8",
      x"e47334e162b9e3d96e26e63aa9ca9e990ac4790d13ed56467a2618f442cd5798",
      x"7a53f4f58668d104a58fc7ec8912204a1aff001bc572c03a020baa17927e6f1c",
      x"41145e18a91f0c3780a637d4ca8cf6d9776d4b0f982194f12ce6882ce887ca53",
      x"18edb534a609cb6b28d294b936118c64a6c4c11dc532994e452e0d7470ce70a7",
      x"4dc65b0cadbf4ef20f43f7c1fef3d5547cfdac9cba1d96644de091f88f402423",
      x"7705293f29c84bc048600ff036b2277040cac9192395b2f9da8c2b7f0634da12",
      x"bde4759f78f1e59fdb5679ce4b7964fcf15aa6bf9a32589178f026c339c31512",
      x"07a91c2875a5605b16ce9feec90df15134d3d620a34d086c5ab1664772762101",
      x"9a5a875689c3ef4b7234a414db2f00e14aaf7af8a5a5db2397f962da84d5b6b0",
      x"7a252d3e014bc05aa647457952bfdbc83d38be09626834bc774da06e815ae7c2",
      x"ac0bc111904be991d5663aa7283a8f8bf4c3cc801e89d495afe130d2362923b6",
      x"5bdd6ec08bcc213c316ea58e74ccab900f4fffecca63d3cd3106f182ee43ea3c",
      x"dcbe6242828be66899d9dabf2648105a3f4e0f5a5174b18b97e5712ae2ba4251",
      x"23bd7716ac6eba2389d1d8a3bee0583d0facf67c16fab30f120a2b03e839c2f2",
      x"67643d11ed6935bcfeeb81bc4af9c0ccdfceaca33328a192d70de00d77f67375",
      x"cfff915066384c71a0c84f73b2aac42c19bf76691b386ef9535adb7a4c851643",
      x"66f43ce5e91f6cd1c3745354e63f70fe0f7868b8130ae6b222dafb2f07b32d36",
      x"912d97a31300a7351fcfca065bc97914cdd25e480b8e4794d93aa7888f4bf82e",
      x"3f8b9c2eb8535913b2c6ab48b7cf7569426742a03914d9dd71d42ba5b56a58fe",
      x"363bf810ac28a6c962503713543b67f977c197caac5c320e167946b0794b46d1",
      x"b6bc2c6f168c99eae742a02f359bd0416105fc4401bdb7e00419c44059f8bab7",
      x"b3595632fa08eece3ba5323753d245f27e98d86ee0e07ba2c6ce4900217b5d39",
      x"a499ef63a57d923e440cd6e1e11220db678c9716d7cabbfb0708bb63d4ae2ccf",
      x"9929bccf3e70a80c781e4b9051ee1d13b2afe6c2d4be26d91f87cc4942df9ce5",
      x"add07b04abc0320fe3b2ec08f13072a7c627cc8c656ef642a561997a7dd20106",
      x"b6aa1e5510a5b2056a2a4771643e7e79f89765bfeb2ea6f94d6844482b22d9bb",
      x"08ed01503f2bec5ff7e3747d209aeb0a2755e98e745e1cef0b8f5bce9cf814be",
      x"d641db74e0671d5b23702ea79e5b911be310f72ae706f57b79f0f06c5664af95",
      x"7c2c6e546d688d4a82414c5bdeadb767c4806de7314de691587b5762afc80cf4",
      x"da592cd429301e046306d0fb9809f6fd599545885ff2ce01b3ee0bdc4a8768d8",
      x"eef8f4f924887c9c320994b3fc85bda82a152bf841a628a81acf8ede66c9f005",
      x"7bcbc8d5828acdfac4e5cf0ae365ca96ff1cfd3fb60438c45b77148b04fab90d",
      x"cc5eec7cede44f6d8fdffd1498055c01c5aef313440bbe334e4c63e530763260",
      x"68e192de5523f7652911d99f07953cd84675ed79053ed5135cf5dc1f66161f3d",
      x"857519c1ca2efa2e62ef1a06a086afb444c55aadbb5b67ffb5acfc409bea9661",
      x"a075b72e3c72d77b013df7ef8559036f4308d9565f33a8d06cf3c7cefa231949",
      x"49bc3544e9ac4587e771c54761eee163ba5e50133985ea782c8f130a69bf265b",
      x"c79b351ac05775c307415966e8cdc9f8f81d4bc144099354e9466c21838887d7",
      x"9db6a1e6b71403ce1781f1090fff69992749bab5250710c1e33e8c1e2549a65f",
      x"339bb0ccb42705d47a7afc4511d801d79975fde25481909e5acfc9e5ff5e34d1",
      x"c370adc8e5399611b37eac092efb744cb4ec99e868a783eef2deb4e2a886d1ad",
      x"e461b93eb08421413939aaaeca2488c0da65fa8997dd94f0fef69f1b0879d7d3",
      x"7f549cb128fc508b13591b7f8ff2464e794433d0b5161723ae678f424e500cb2",
      x"fd721a7021a103dbc7ad63c49f2d994e4c19fa1f2f6244e6d6aa61867ffaf2d5",
      x"384afbaf1d9b5d7205622a53ad16b80a43cd424a90fdb7e780cba129bd7263a5",
      x"6b0530ddcab5e8bf794bbf867efa87f2ee0465c8607bf14a30fcaa8d73ec212a",
      x"aa030f297791899fe351f66ba827436522590a060e01146f479b395b112fe319",
      x"a897f88e305cf7be69f0c3721b9075e840c6ef9c7c32dad17a3804dddf364340",
      x"e60bcc2616f62e7fd7be5c75b326a2689a53935aad2e6f7ae1edc7a9382ab7fb",
      x"765497cdaaf96a5737757dd134d23587603373039d9ad574bfdcfca20b02d92b",
      x"847f4ef623771bf82844fd7cefc6ca28b65accb50981078c6840c62f64b70ff0",
      x"b725708a5ba4fe89e1669cce41cdf6a63b2f269aea3e97efe9e140e576cde89c",
      x"13de00ac82d662e73662562a9f109097c74012bc3f4e167d24ee1523ba8d85bd",
      x"a4ffcc511619e938cfa6be1b65e91476b1260c6333e18d0367bfcefbc7854fae",
      x"fb186fa17cd98e43f7acae18eb83af3ab0d97566cac5a368e6ac317b5677a026"
    ),
    (
      x"0f35196d5fb9a25c59f132f9870f2588ec14cffa3d8ecdc339240aadea2e6199",
      x"6affa2ef1d57111256597882842013a216fe4a54feb5b1b30d23d85d58f4d585",
      x"f00812655c47cef2290142ae5b4ca1b066f2d66ef1c5228a60ae4b20bfed4b8e",
      x"6b09cb0ccadcb8a32b9c030fd3f74d494e732bba54590cc82a18f1cd21bbf443",
      x"49a0864aba8ff5954d63dace230dade7b6a8fe5cd1a3813f61a535418dac388e",
      x"bd9a81be515049fea42fa3c690e7b0752173819f882f49fc3abc9cee6580cffe",
      x"1512e5d625a2ac9a5638227e65f1e7e9fb42cb22c3449901b17f0e45b31fa5f4",
      x"6eac9e647a386e86850d9f4564e52a333bf5252f66972f559000115bdcbc3b6d",
      x"ae1f37233ddecf95da1ef5255d1a37c1a915140b9d3aceaac6d5a7dab5a99e64",
      x"0e02d1ab02cafed571365620393e5c1195316d6bc41e7d066c9390bfbe1b9cad",
      x"9ecc16196c9ec084f9c23ca409b33b6402135ab4c524bb25a55a9127b9503b3b",
      x"2b2ac7768b0bcb4360bd5a13303d306142b8e8aa8c4129905edf6845cd8b1ddc",
      x"85b45ef6c68d6bd3cf615e04d1c781e52ff98602ad6b6a2954b825e0ab79c614",
      x"94f9f3852649d1ac37ced7becdc0dc3b2369917c084cb5dcae35a3e4fa87eb3a",
      x"9b1e8fbcfb0a6393598e70c6497bac57c9cb5f65a7f56e1a25b3a9f7c7c981cc",
      x"e6b7a552dadf82610f5989cb89d87f683a344948bb5c6eee6d011c0d79cf7261",
      x"1281b20f156cad3114e7310498bf5645b8d846913faf50ef4187cbc4b60aacf4",
      x"02b45dee5cf83676946f81c9387b399533ac42cd0b4557b7e6499aafafc1160e",
      x"511829641642896dc58b16de64a66ec23074972982898e4218a09e09adb7bede",
      x"478d009328a9fdb219b6c63f28e43b951d337aa34ef632b3b341f1894133782d",
      x"d38e63507139da648588187b8a3ed8fb1a09f4dab01346d995aeac686f0dff5b",
      x"46de4422c0b14f756fd238a1b843717cee078ce2c7ed165fe245fcd96f34d8ce",
      x"ba914419cd8fba0e743aada3ab31ed68c87889e25cf659981a2391101ba9fd47",
      x"5f46ea845831a4e2319009593aa728bffc8775df468d3310dc97ab0170bb280e",
      x"7623fbfaaebb5797cf0dd06fa64888153e17af0b4b5f460e394fb39714bd7571",
      x"123223f9f6493aecd44d2a7c3580a3b54a439c7a8075fee0ddeb9a4b0a27dea0",
      x"0373174996a285a2d84980b33b5917438c57cef5dbc61e6d376ba1d1524fb397",
      x"14c386f5b8148f16acd97e15979e393e7f3973db7900fec7533f4e4e84693e1f",
      x"26769989c6e5909294f9894c328919631dc44255e4cb224fd3ce5ccef7ccccf0",
      x"52618eed9d8663147bfcdb4d06464e5f93cbdd6dcd3d10decddff98fcd9310bd",
      x"9db1028ec1573173d0b0a1a3180734f1afc701a3eb09efa38afe7fa9db2be611",
      x"07cc147a0fc43b0c8fe47e37118ad4c63a68015549e2406a3427cb42fcd4f4c6",
      x"957e43780798935526d8f38d970185c95dd0c3d09a9df97204474e1f53ef2544",
      x"48b659549e08ca9bbd3c120d3378e286299cf26587aeaea69f36efc4422d4e0d",
      x"7abbd7fb6331b135e6d8f8ab568c3e2cd18a90c03375e7469c29f2cb6bbc59e8",
      x"7763aad57476d7aa1617dd6b338b7207c3fbaa8f053def801ddb080f3acf5b41",
      x"651908aea8fdb5b73c86d6ed5b7ab2f386e541b47ac790abf6188b5616cfcdae",
      x"c501ca97f080ad51c9da4bf4266f99761a4663ec02c9f54dad4af75096f77e1a",
      x"0ca893f8619cfc1b8325afcad25080603809a12cea96c6cba2e19a5595851c5d",
      x"723161768d2b1cf48452273f75cb5bb204f440c26ac955d341d09696558f1271",
      x"bb5f89d3969a50c76323dafca21608831d1d75f8bed78956f45db416422f279d",
      x"323be7a437ffd226c99ad8d43817217db505c7580b00abd5d0a68e20641eff99",
      x"ea2f427d18173c8a76a82c425b050226ad3a56acedfa3a97342e7eb4e9e4edd1",
      x"56771e82e7c1206462970f50cb068110aa9580396e709b8a486e9b394b527f41",
      x"5c6c8abf4e0eaa1a54941a91c84b7bac2a1822d3b0e92f383124a43e039fbb39",
      x"9d3d8725ae0d6a66bab03f2d8a45b5b2f243e77b56ee7f68812c9150d7b0c8b5",
      x"b644e0bd4902bb81f6bf79412ee188d4eba9d66fcc8e570a188b1472b393645c",
      x"b53927741bd792e619d8f6ac636331400c8e047bbf629467d0b4fc4034750f71",
      x"e74aa6b3714a549d900e9ac59830ce2421813003aab175e4861059a410f2e49b",
      x"33b4e825a65545c13d393c6db565e5ae082c2ba4cfbae709c8223bce03919d36",
      x"a5f8f37c3e4c1dc887fe09796792367584774ac7cdb3e27d9ae7b315da9b49f6",
      x"437a93bfdf9dcb60efee843a226944ac8a23495811101921c093458d9d57b219",
      x"77c0ca8da10f31ca4926cc2b426d78b03b610754698a3cde5c28ee0005f5f502",
      x"46bd75832625b428a77119bb282467895f80a825f44d5ee8165e717c70f2c731",
      x"911abe0327423ffa4c570be29e90d5cf368087d02ffacb89cfdc9365a1226773",
      x"aee86cd46d02c3e371180697c1f43adafeedbb176b482f78a692bff1ac51dcf9",
      x"49e9adedc84ed8b8efc1555a7e4fe4e1f5c81decfe2162a393b0750ec0f4013c",
      x"25c0828ed6c6c3ee35fae87939c0ce953a6f3e6e286ce0e93f8aa9ced28bfbf2",
      x"65ef1947487c54329195eabf6cfeebc936c37e0f0a343b546f5f374e63d1876d",
      x"3be412769465ecda27ef91b3025679a8ac8cfdaeae1a5b7390462fac34d72bad",
      x"5f22eb0fa53dcd3273194fb1cbb8e86ea975898fe799567753e533156c38a602",
      x"d57440149bdfc22cf9da794e3a385b74298288f79fb8a7d0c2e0f0c1b8cc1999",
      x"1e1bc41ff557d1add311a3c707f936edfc3d246c00fc3ef89361f6723d12dd83",
      x"c3d5b39930a7e2fe2bdc7d0ba1292ad9a92d542a5f703da029c97378761e7792",
      x"b93089e360b6b573f919aef78584d0fb085ed2df86c8262cf15cc7dd51a10b0a",
      x"fa31f1aa5a2ea2a78a7ae01b256ec1d63e86e2e39792bdef90cee8f58e97b882",
      x"d92d2657c1b551cc3b3bdf6313e81ccf0be74f89571d3d7e80fb028ab08f2c09",
      x"68854e35d623012e925f5c90e2578a9d7f7005aa27cc07057f94afb73b0b62ea",
      x"fd163140edd999e77bcef3940caf1548282006c6c632d2bb8feb1569a51ee531",
      x"e13dd84a6f25f9c9aabf6af6b0266dfc55e4fb574f0673897c264477f52433ce",
      x"5ee68f0229c288a5ba7454e86396a8275586a91cb62990b71be738a58580c966",
      x"bb65e596d983c6d88d03f3f26a80fd98af6d2deefbb2da5472e95fc42a722aee",
      x"43db63a047f459308198b7ad263d5e172e46131288d6709be4ad68fadb5ed4c4",
      x"88b0ae23197744f31ba9e3202c98da39d6ff786c87be639eab159577917d0c02",
      x"39703554caf11eb8f60db4cd6ddcfeb35e45b9061967365db62cb02fbe0c60d9",
      x"bf5024392e47aa1036ff18f875635487cd633c3068cf59ffee2d289e8dfe86b0",
      x"de2059a941cea20629d8803f33ba67eff8eee57d70a78f9617bfa8f37d22edad",
      x"77a3f857b714fbb0c32bb6566f101a408c5ad5c765da702ccb4c4b9cf58dc052",
      x"b356e45b4b08a62f09581e1c7a17a151e8d20a8e573e0735c65523fe5cfb2c1c",
      x"8f1026cb0e71d9110fdc1577d6ef36186edff42d9346349d93a094be091ab7e7",
      x"0a1cb2255efaf027b0a09dffe4359e8de43ed07caf01f76e5c4c8160bb0ed208",
      x"d9560c2f3ee950a5fe66d544ac5d383e97606ee429ced588e480ecfdec02bf86",
      x"6c673bd9a58857da5d9045e08405ea06437ef6d3977ce13e2526c81242cd1e46",
      x"1ad7e2e70462e2046e10b6ed019c76c5165e4129ba3e2c5d58eddd6c6d820296",
      x"672b5f1809632454db9ffb2934e7503b32222fe22d81f0cc8681a7dbb49cff67",
      x"f55ea31dd4ff2a2de46afb0baceeb56ef9529ddc53e20945fcc6a675ba342b8a",
      x"2df6819350947ebbcefb3301a671d6d617919cbf9c9e420a4eba02393643aa79",
      x"fc99458407a4c7abe5c5a7d764b2b5648a6553f4d2cb11d16d9bd3be79f3538f",
      x"88e622714fb33b68c98c8aa58b7298c075501fd37bc6956c4f281ed30287fc95",
      x"37ba738c610909750adad21e56e4fdd68340eb63464b416218039068906858af",
      x"c706dcb4b03c5e9bc1db321ce4ac4f04a4ee0a9e620a778c4e2d2177fc738f12",
      x"b7c7ce43df9acbcfb04e169ad62e6e760768900d341e5faf056a2dd57875b8bf",
      x"0cd1c293881379b40fe074e0c2158e9271bd1fce89498b39359c08a66cc73391",
      x"43d1f9ca945179d5f5c96105cbf9204cc00231f57cf283329ba6a88d8c22ccaa",
      x"1aa19cdbe91aa858a439e6efff3e764c32a3109e51c530f97310f5f8985019f5",
      x"0019845e141fcb786d074fae12004dee772f3cf98526fb8fddf8f3a71d098ff0",
      x"3f206250592d4f62199f27fe06ee35e98f2b7fa915ac94b5223e0d5e9197cc3d",
      x"a57af98f14b5730dd609f5431889c90a995bca06d431ca7fadeadb781650ab88",
      x"f4fb27bfd57245c3c0f724704df77e712b4aa217a07be707d22487818965d6b4",
      x"67a8e59fdcb9c0c96f30e8f474d1408f180de0a19b30c62db8a8a4fdb8910550",
      x"fa9cd5b43c4613e88de84f0263790ecd3b353896dba2e66e3908477304a2b025",
      x"4fd21adf6880d5aec11b2a58f281353dc0b56803ac71b70973fc5ffb1bd06657",
      x"aae62eea0ab041ee4ff4b1e6b5a6ea3c9653c1462463e621465b86153f74bac6",
      x"a4c606411a098b48a55471ae577f35d8654832b79830876bd601af87870d0947",
      x"aa5a8ea20e17390ef7d8326250a27531e5b5ab743bd3e89385a1ae9c4ce7a6ad",
      x"b0393aadaffde59493ad95383baed3a61719ad15bebde7a6d7c48af6a557b7a7",
      x"4fedfa1f66924fafbdcd56f5b843bc4e6ab8bc3300def2d41457fa37a89a4a0f",
      x"cd30b1c0d8ffceeef69d1967d60ac636414e72b4e11a240bee76081577a5d025",
      x"4301845791a4480ecab11aabd4467b7807dfe6bdabfad6ac9051331722f9e173",
      x"a380a76c57d260eccd099cae5f7d3528b1a83c49acc5d75641d01373d2439a6a",
      x"a025abf4c751c4f4d115df886cb1f6196b79e892c98d059e81127fabdd0305f0",
      x"470b0fb82c81a488eeabd77759e7309257666e71ebee82dd78bb94a6a3c67bdd",
      x"d6ceee9988c4d7d3823dc023137b087c3143beb28768be29c8d8b5d09bbc7860",
      x"794859f097a1985992c9d6970747885c393a25dd3b717970a0ea61e17943fab6",
      x"cc2dc74cfca0b40927444077fa57a94a72d14500a8e2bdbfdfe78e7a7272ccd8",
      x"61f6e509a08ed92f5ffb7ccfbd2e1ac2af01802de00ab7d6c339c3cb27ff3da6",
      x"bb5690ae0b47d8e8740af6b38ec21e29ee6358d56de01bf057306a52ae43185c",
      x"db25af42b305a8dd33260065f6a1d793428fca361c489e7523156ff6ea136200",
      x"9b8092cd8bb93ab83a96010dc9d6dd4d4631c599a69546851059f6add62223fd",
      x"8d53826a7ab157d3fba416d71f0dbc3bffda52478acf82c7d7ed56f8665186bb",
      x"9854a73862987ae922fe61b44f66b624d73a9e999a24474750524dda5bfd79f6",
      x"7b4ed1f7675bf49873fcc619a5670a3100c3edde7328b03cc30270f86fda0d7d",
      x"7b929b29575aecc623ed17b8eddcf54d31519e15ee28cbe08a92038e43b18a68",
      x"3a94933d30d0905c75046140e17a454349cc09aba492227af2675272dc4bc0c2",
      x"d607dfdaf54b24c5db2a0a8d7d5715c68342c6e624405409c25f4b0b98b4e19f",
      x"1ef5d3c4569c37109f020fbb238b5a384fb2e5b088f7a2156c8bcb14e64152fe",
      x"38a0317ef27eb47dbf90082d0c97226cda90dd9e9f1c219a03efd02f16cd829a",
      x"3f1ae47a81b889091d8bcb575d0bc16e05a24adf03b3b2b2f7d09464e8344052",
      x"b097f1444b459d0c52c8047e9113f9c5df6972df9a513e15b9599025243d8ac9",
      x"5f46377e1beb92b22801059a943424cb1b32abb818938f18d08d156a5de36968",
      x"27261dd89fa7c52f18011b5ac095b7c18650278395170de5b74b505d30ba0ce4",
      x"9c71c6ef2eb71527248a9487c02905afd1a879931ce75781be0a713451d010bd",
      x"363e5cacc4bbc5584a2c9d7a269638a7618b5685739cb5e9063ca4601e5dad7e",
      x"817612dc9b7f5dfda50dfb49fbede5aa99941217266c1701111cbbf312c20494",
      x"0eae0e11d553213bc2c8b3e5ae1fb4627002e68f78790834c6126502c175756a",
      x"0c1f238cab4a280d4305d2fea360ea1ce2b449f4ea941109f27712309c52b7cb",
      x"73194da1904813629c6b9726582b3a9e971eb1de2cedcf1f77f9da3c75efc017",
      x"f1025d961bdc6cb94a5f3472e4c6cc6a7c68d726da27ab40f3fe824409de39dc",
      x"00aa6c2f2021cc8ea06501469fd583df5d8d74f590c49eaf17a012537d411af8",
      x"97f36c7b223023c833e3c29a909a59c3b6acf358349ac57ddb6e4cbec719767e",
      x"37adff0a48bc2558a83dd924037765e297484ecfb5bf15446da97dfe78419e32",
      x"d0c77de25b9c327b8e4a4936093812517d9546324fd2e64b322b101ebfc1c993",
      x"15cd146e07f509c31da07be010d833fa16262e827b93a02cfa816896cf6c4a68",
      x"77a18f8a5488a2d171378247e854bf5e6ebe4eceb29d5a855174324bd4f56b9a",
      x"aa373684c88ab32518c4305e2a6a00aa36651a7b4240de691503a68502605299",
      x"c232d33b0ce0f248ef02bf6c486cdff6f6c41fc300d20fabf509eb6bf76e1caa",
      x"fde28e641d21c08efb0520e60d9454255f8a4141cb3cde2dc4ef5da54e50ab7a",
      x"bce3a418e93b090eda5c595468d21a98e96d055ead86051d3f2254bdc3235e7d",
      x"fbe9fecc94b2d9ce914561bc350cefe4b420550ea4a918f4bf9c2e54f4831012",
      x"0a9928b8f8e9cb9a07e10f9216275255d9cbfb86183f773d2b4b78781d241e89",
      x"5e83544d610c300033e04a225ae8f2ad97c04db1c877c0aef595ae08353cd0aa",
      x"d06511101ed640c36f6b56818c4f985f1cb0bbea62477aef9ecac7bb0c485280",
      x"47cdca5ed468675cf887451bd38ec409fa020e68bab61f9ea3275406de8cf6bd",
      x"61d5acca3e45db2751ada3daa5083ea6194e28beedc7a036e2c5c780882c229e",
      x"d95710cfc77a1c09ded98dc1d2e9a508d2fcd9d092d6abd273b286c0cbf1b68f",
      x"7e03ee7b0562e2ad3c118f41455a0f3d6a2ca03f1f23a22f16c281bcdae42dc4",
      x"1725c1a0a3d27bedaca7169cd6af9c7d5bfded4688189e1c12a11148062c947f",
      x"0766cfd3085614e2b5d14177a6177a26cff37c79bc51c7cfed18f66eb9d73656",
      x"14c4170a9cb6399f2ed65627a82cb4097c7548712bdfd181dfac35b3465edc1a",
      x"7bd4c432a64ebc901cb22c9496126eda3ac77cb927caf3717cd243a3478ce4c0",
      x"bab580b97ce4c32a62ac97df087ba49eee7c687ded1b96c79e290ed252e4cb35",
      x"61c36aa5dc674dd47340bd2653c293fa0ae316cf1a7490f297053b9ac74a051f",
      x"d95a85d38955273bfb5d1b53407b8457faee8d7b83a138cc08d7e9d9df2983db",
      x"16a7be8e691eee6cfe67b7be986faaf9a6aa5652177c43b0f2e4f23f5e5e4d15",
      x"5e420a7f9430caab70da6cc45bdea23262fbadaf872cf56f4425e8d19959cc58",
      x"91e573db05c8e773bc897b93e5ba75c1156077454e91699a55de007a3307a634",
      x"3b978cb85e0bf9ba799f2ba91c314ced98dd911d114257e5080602397e9815a6",
      x"0e3ddd85b5c7af87592246057f00e501bc4dbd313d0b73c63a01dbdd0cb59475",
      x"fca6b3d9c7a79d63505ad53ca7fe3cedd35f98cb87242254449e5df94b62d175",
      x"78316c9ba105a20bc6d6673c37f062c6c2ff51374f891b2b2c0a626bbed37f7b",
      x"24774c1f0d9add296511d37ae8f7cbcb707200efbb2876d9c7587956b0eb3291",
      x"de40fc236005d31c43475fcbe3615cd042a218f6a8a3055b2fd9d2d64d8f3cb2",
      x"d8a678f12d8d3f2a17a89a435de13181577624ea7bfdd7e88462b1c891eda8ee",
      x"b85a3f5dd26aeade617d314bf13006981cecd17ee483bf42919c32a307536f92",
      x"b9b7e98383c0b64aa0b0c35fbcd950a51023512f8b930806ae75d0dc74556ae6",
      x"c2ec06230cf8b8db78feba61a843e49adf1a8020a8373bb51a2246a9624adaff",
      x"29ab7855b487e7923546212dcd772a6654a8cc73e874b3919f62697e18b928dd",
      x"b9d506900321a75612649d9c2b28cd64027b9946daa6f0264ff7cac4b31f277f",
      x"91ce2ca4dfe27290595c696b1062be9b03ffeda1b4e9715a040e5ed5ed2a1fda",
      x"70379e1a322c27f5382389e428424f6c2459cacde4966804b78daa42e2ed31e1",
      x"d8abf50d855d03fe1538ce0d31e45d7977d60f5b7dd4b0c71276b5e6571b24fe",
      x"26a36a21f24feb2f27e922ded69495b3ef1e633cc051bee431564deb7192aeff",
      x"bea981af1111f93744164c2cf66841193b30f4f67e4a42f6385986e6d2714ee8",
      x"3d3227c5e3ecbbcb2a410083b64472d14692f9295020725738f155a5175a8669",
      x"e46bfc8736d58df404183ee555636c937ab112b7a2d779e72db9beaaec2dd722",
      x"f972fe1c11bb1844f624b314a78eca472d280856d8b4d92903bdb3513d745523",
      x"54e4460688ea3af26c430f84aa1b3182290c2173250246834ae3e1310bbf7e6b",
      x"de161e7e38d61ef3b0b736eba7079d2a49c33244644ae4a7a1d56746c8bc3f23",
      x"978c4a9dfcd66a93262fc525c82c0078da0f8584a48bee7a9f750cdb1baa7de6",
      x"a6045cd9f11a99586e36996267428ba58bc8ea45c684b7de14d0b985e643e490",
      x"150f3b0839bfea53f80c82aa7207602dc5fb6d7cc1d8b8abba18ecf4ce81c399",
      x"1a3178c6fc6da731e4dff074dd035be7142fa6ab9072f2071cd74e5702c4bdc2",
      x"6d398f7e47afdde10dfa51cf4053861ce8d0df2150d868176184a850b5354460",
      x"7736bfc84d64a41d87e0a990c7e571301507ac3f02a15fc95795d16295aaeab3",
      x"626329aa2b0d907ae4703e64ffd7ea8d73698e2d4a0bcb171d9152a1dba499b1",
      x"b7996d832a9fd90f4fc8b2b9a657d009ecb1ad9b5057412923b70520f0d95eba",
      x"9d5ca22dcb54eac87a038caf3f89cd0d5cc59a4ac383055dfbe6c3ed61abcd55",
      x"05abe402502d3752d96209f53056f92be14a8f913acb060896f8f7eb1867c0ce",
      x"6c5d1e6e0079b72ac9f8349c2b26384077ab9c1e9b1776a979cef50fe92af716",
      x"300db04ded654309b298000ef7a39a6ff40a34a1a449dd7988e686dbbf5af75d",
      x"d9dc89efa483453bc887fd631e470df012096c072e1e63ded901166a1d1a17eb",
      x"77ab3004f4733b30edc9f87bb0f89be37bcde5d7bc624f9945b28aa32f96d498",
      x"596e1db17e6f153b92d50be6d32e101595b58200bcccb72ab56883a67669a9ff",
      x"5b5f3a5ea4a44d6a0e7ca1846516d1b65f601525c023cd4e2d3eafde28d3dd51",
      x"e6fd30667316b6fc6c555204198e80e1ee64a7e148b8feee867761485f64b63a",
      x"5dd2a432bb1a68a11c2eb845af244f9858e5da1ac4a231234ec2de5404f70917",
      x"15a6df6a970752f0da469658b1ef434cc49488bc5e60049532738828505e4bbb",
      x"dba26b59273dc2f023fd4c45b325b06cdfdc635ef5cc39dc61b29d9a97fd99c4",
      x"793ece13776157bf07c59a40904e759042f6530d9e23e252e6f0a65ffca71894",
      x"65c42984e1e19bf74a2333e24830908ef7476cebe44bb870c7621b10d546e3b3",
      x"5dd1f559ed29ef179f48352b40b48a9450a68cfd52a9eb9bebdc4bfdc5749701",
      x"20222e6477d82b3b75fa202d08212ba29e923f8f30066b378e3e0aa6226c626a",
      x"ad8525763ad11defd11ce6087e029e948facb95f3aa0aad9566af9447de2b8d7",
      x"f02982d1c3571280682ce485b318a61e86ecd6f1688017ac2d2e2139e6c7d644",
      x"c4a21d6ec825a9410d1046ab78e88f51ba9dc2580b211436d4c91603fb016706",
      x"97b39777faa69438205636b3c1ac9b3b4382e468cfe40a16dae5ded7f0e9c6ba",
      x"8e28c27c3af8fb99839d57cf75818aff509f15c4a65d61757c092d649b0de192",
      x"5fd085a72ccacf965936b7541dbeab92ca579089875a304c911ae5345e2d4e77",
      x"d3bcc63335f660f7e0ad8751118c9ee4ee02e4b26d2ed1dbb58e62a4974532d0",
      x"2ce74bbe44ef20d71d9abd3215974ab4193e06e43fd462f5faa7af76cc7944b2",
      x"f577d21aef5db006e543a4cf8d7026b685eb1a5f70644326854cd7a7e06cfd53",
      x"1629dda0a965a9eec59629d60d0eeae66bf5456de8c51277595eb7d1a70ad3c0",
      x"b710572037259e9d75634ac44229135ed6ae4e9518dd1b85b3c72c92a677f12d",
      x"2d8f05e16de9f1b11be641d62a63859e152860b28cc1a89122dd002d3102cc69",
      x"c0519a5199a04d23eff45cf4c7e57969d3fe191d28f39798681b2ca1dac5ebe6",
      x"feda391d279202f485a8790fa7b85a9f7081d299c60b456998fa731fa0f72de1",
      x"2bf7a281f22f05415222c9bf3e7b5bf9fe7cfe17cb89d1ee2d4109244c10bed6",
      x"adddbe7182badd7344bce60d1213b510fee100f1d012e1d34299cceb9ac0b64c",
      x"0e4af6dc0d415b699b277e05133d69bf9590cb6d6b6352564b0549913ac45fdb",
      x"22e17571e043a16acad2b377a5db06472905a9e9601cff73de848a8d82c7fcc8",
      x"a566ffe7fd829c50f77df8ca062ecddf24b968f27bc1c43076ee5f876f636887",
      x"1f0a3937f10e5dcd674f81a12096c7d609c94d2f98ee797d43e99bada115fd5d",
      x"7408f78bdf2cf6791c29c2f4e753e07b98c7a942b128753e7f9dc6707027933f",
      x"ff6ede2fec29b029bdbb17c24e58aadaa3b8fa2016206d760ddbeb785a744c69",
      x"6d494e78ac432edfe27ab6f03347adaf680bfd964d8418cd98876de980914520",
      x"ad4ec5ef8aba2b6408d41d036d80327fc746f12433155c237a2d9354d871b68a",
      x"5eff5f4025d614bd67a547361bff5fc96326877ef518b07bd47d7d9efa0342a4",
      x"7291f276b09401add332dbfaf48cb6fd4a5da44559fa2caf8b430284e265452c",
      x"84f3d1aa304fcb3086ad455f9202a3aa257bbd8076a9fb654e49f23d1b3b3b82",
      x"96c869e3b082adf7e71ec526aadb6a26d32bbfc216a7bd2da2b6350a342d9fac",
      x"70db8bd3266b935b43406ab627dbe3a4406ffa7c0d78e9de9868761f14dd6e40",
      x"63b1fbfa9af92c7e4f3b7814ab40b9b6007898452f80d02db91b3a24462aad20",
      x"96affc64bc4c3c1072e2f08604b2743816f31a1d34c2adbce6862effae52681b",
      x"38f91e521544627aa681d80d09d7b321a9c01d9f256276c53d79505c94b6b5c2",
      x"8a74085c589f95aa2a92a9d7ca0822f832d8b6d91fee769da95508900a801e25",
      x"0b5b156944dd05504010bd4e8e3756233836576286cc9ffe8f8ac7d76abc5e45",
      x"eec11d7e759bb43a27560177cb9be2bae0ed21551fbebc71fe9a88a2ec1dc8ce",
      x"8bf7fca2366793ffb9af482d4a63add17f913016f12b835ed8b2e8aee195234d",
      x"397a6451b4b336f712d956f3297a436c48bf9a6b20444ec09091c17fdf71a4f1",
      x"60a4a7c9ba9977baa1bdabdd25bdabdc0d0a3a6caee5086f7356b49745209ec7",
      x"4bc7a597e4299d0ebe41a54b916b6335752345e307f91c3e18045cadf8ab7368",
      x"c45eced401b34015095e218ace06eee9f148b12398d54b30fd301579fbae617a",
      x"96059346e7465afacb140003ae518d53bd40a520f077e14f4453827250a65bc9",
      x"cd8c4070fac8c3fcba04bf71dc1abf59bf57bb0a09fc76216297230e5baf2158",
      x"5b1ec48c8dca9dc4acdd6566af338691d39dbd8a4213a80b6ea57aef071d0d63",
      x"f99d6e05472abc53d74e0c5f4d03198a69d4bfe8fa1d8461ef6d927b269e7cf2"
    ),
    (
      x"7c1ed91d5125698c93e22681983da5529445b3d16d39698947ccfc43950f9456",
      x"eacfbe7b8f4d0c60b518dfff74fc4089fcc468e3986a92f31109b0cd3f68247f",
      x"bcde88056813050a24b7b0b394764f031131e8b6f4abe7279c296c967fcdb060",
      x"67e8640af2000229a2d0683f7663c18e7a4fbf210efdb502685f1d3e7b6d9834",
      x"00b1821ff01381cd11b23ac4cf13dfdcb044c90530cb94822ee162e56ba881df",
      x"233fa7e3c1dc0794667b914d6ab1f07ca6ec981d0155050ac7c36dbd5d2eceba",
      x"b70415506cb79c88883b060b3eb334e8f2d193f43d83c3a06e33204373f3d9ce",
      x"84ebe595a9dd7aea21b3664ca308b92d4affc9c389ab3174e0b106b7f37a5480",
      x"f675cc2f8734b2a623e78bca189f38f0c03b1bd869c05ed8aee276703d8c5c8e",
      x"f5f77e699ff80f4f087e9ee892556963d86af41c6b2be7bb42ab85035d17d4c0",
      x"a872a4a96a38dcb42197f470b6602b2076b480a01c5aeabbb040f1c4957ef901",
      x"5c3be324a9fc04c4409914d548901f1780f9263a97564d96160c05c07975e367",
      x"dd7e1142eef3d617ce79f6a55126a766223c16477ca79a5da8ac83ec2f9c59e2",
      x"e13aa45bda40cb9c6fcdc62da2c7d80d4494110a0ceb9268e54fad33362811fe",
      x"fee10e926491c3e4a200ab20f3491f5a573e9d28c355a2b60ad6f7fe2202af98",
      x"72aabfefd61ca20b8591bebab88c7b8d9b1267e0c0358787c2d0dfd0486825d5",
      x"e1c093d1153ee21a21c82c4faed3a0f403529ac3b055e7cbfe49a027dcca594b",
      x"9fa633d77d8e9c100bbd657cb6458a7ea2a8e34b30546101bbfbadad9c42e59a",
      x"78a1c3338dadbf56c3b015d4c1362e38d0b589fceed9134cc82a1bb55aec5f79",
      x"a30e0b3c38f2240a49a8aadfbe130683d555367656ed7882303d08bd5cc55723",
      x"95f2397de2c08499a0d10338c718ac314e5c1b952a22dcf11ea1de65916055e1",
      x"3470662ae307fb1e8924474b99ded6c128b325376789afb100805bf993f1fd10",
      x"792d1a3d612d1ac78850a3a9a4b4ecfe41715e2c228595bfbf6cf68bd1864dee",
      x"153cfd6eba3a57f86f1fb7d95c696dab745c0df034dfaa58e349b47045036373",
      x"cdfbeda281d3cd136fe5ea9561cc819e77491888cc2f25342fc5654e6c8ac4f9",
      x"fe107916f5168ab7bf4329cccc289af22f0c3bc1ed66292175c251a81c063ed2",
      x"31d3e75d0d3a6d979a0cae7caae6d215d32e1b23e63203ff3fae8d57276f737c",
      x"c734621defb15da7299b7b68d2a9efa080210dbb664d5886bce0657c627182ed",
      x"344b1ffbead30c0c5f3f2ae57e468969768dc3eefb39263428e78c06969ac343",
      x"7836a4f5c542bb503e3fa3bd8bc5d9a9f322a75728d5248d9405983d1e476c9b",
      x"535853e8b2fde9ab34573e98c5321f24471ffa73bf169ec63c4e4eac7d630bea",
      x"1a67362a4534777186a757b87353bcda0d67b5ba23b1e647db28c2875bfd1414",
      x"4b613e95a0e5bdc840e0e7da839614a50dfad15d8a0fb5174d791239b959212d",
      x"5cde6f281ede15d3a86ce3422d17438aa5d915583874740f6fee24235c991edc",
      x"32b05269b761712a5234414b889c516556cddbb4f73c84abf7cb46262818b77a",
      x"d7496f285581927f87901f884650df59416e728b782149afdb7471550b63615c",
      x"e664f60fdb33a2f8862367b972d1c22b2a3be5b36a06a52a7f195af547fe08c2",
      x"ee0a3e01a9966a61845c6357964ad5c575c8702be381cf30ae4d246e0f79a3fa",
      x"0b0fec257db5a2f05e13ea2a1ff46df6115cbd1dc0f84edc50a6b9508a5451ab",
      x"f1fb951395f33bd13aba2ff4efbe81409dff89ab09080515de72751aef6bf7ac",
      x"7def097e09d1646c0d67906e26f3d283be855074691a8277eb5e76d2eeb41188",
      x"75f43499ca9b1e9d8763472e301bdec001c0075bb56b15acbc404e70fe27b040",
      x"54ae50f6467ebb69b71f5685012d9c22f1da2779a79f2b6005e3f9b80397d3fd",
      x"7597f21624f1af74146727fd8204c0bf756d089f27023a48e0c8ac82f6de3b2d",
      x"58ef6d58695e0784077d1f1ede65675f2d275f905b939d5d7d2d3521a6cdfe50",
      x"caa50a5f5f2df0f677e216acc89866595f8643ab9e48bbe3c8beacc63e6c017a",
      x"a4be4ca2c7364f024920be8456765972c64444f5791e6fd94cff26eba919c53f",
      x"d663ed8d7a0af78c1aeab4c55a19f9c78e3b510b3c87636b46ca821e648aa7c1",
      x"ec93f1d83d785055fc8213d2d0b84dea82a6c6b609d371635d11f562a96f650d",
      x"2698d19303c5c25ad679b20de6c9df9e98e5435fe09f4813fe16522dcf5b0553",
      x"2e3ddeaae207d20ca1b03e034e3f99957a0c258e0b32771eb480605b3c35bb8a",
      x"fd16aacb7de13d551919c01f25881861c6bd84191ff3fddccee3dd19ef165719",
      x"930fa10d8c096a30f955ca26849780f5e8081b20122857582aa10f025bcd06e7",
      x"ff619c19e3fc7e3976ffec4606b8a2d276bac4277639a7eb8994da478fa6a51f",
      x"7bd88d8140dd9f11353d83ece73bdfbfba04aa6d19568b4b58751fa57834cf2d",
      x"f18107736c582c2cb1ebeb9bdbadc7d6e56b261fe15d70ad2ca8148140c6c798",
      x"cbdf5e309c9e7a282405746706d2a3c5a6aa97e4a9a57992aff863a1f8204fb0",
      x"3738314b1aef84d10e1cee1ddee91b64ee968e361413722dbb73bb10abac403c",
      x"606e997a79056b18f03a4a8e2f330b4b2f6c63906048b0be3faba5bc85529ce3",
      x"a70fe62727ed5459390654e8ce57bfd6e7b5ee59710b8d92a084e5d33d9256ea",
      x"afab5d26b053c5c38a1dbff5359020529beb874f868766b77885cce77a262c9e",
      x"80c46d1f136a4dd3edcf872125f647e389b98a4fdccb9c1de25ac6730bfcf57e",
      x"a74e98b9fa58d543c3afd626a9974d8dac2d42b30890101ad8b7f8ab2079b208",
      x"98965be0e587e9fd8c66c999fc078814c5d173cf6540a9e7ec4800f435a27a5a",
      x"7651890a371931737c467028c669f83ee8b2169f8c87887c7d26f2e2811f3b40",
      x"2e8208513accb1074fe6a541a71ac94f6f7a4597b12ffecb316db9750b955e32",
      x"b85379790d31a418e654c8f4bb036c5d284a78b08c89c5b7f8d1efdd5f2e818a",
      x"0e202a37e786790ffc95cfbe1a9e08e965ef513761e19fd384bf64781f4e2c06",
      x"67c1fb2a2220f51492e45601caafce4ee02d1365c7bcb9d3cd32e8c41715ce4a",
      x"8db72d2d32aa9ad6b4215fd6f9c230516ae60e8c588b6cf9ab479c1509313e25",
      x"dfa8ee30f8d819cf0710f6673388beb87f9983f099a148b3e2c9d061b0332141",
      x"c2968e1ac5aa578eb17bf4a37a1cb553312868577b90c2e7a9db17a25e83f272",
      x"8337b2e3a81792ae4f906a5f9c74f2b8fb5cbfc0858385360157478c1b5d7427",
      x"9e368ee8c4afe5d5c536df96daec5888cf9249b1044688b2de07d17bc5702144",
      x"fe444a2ca4dfc7ef6bf9e00d20d9f72c95e30b3eb7a10e8d8f4fedcb42d3571b",
      x"0a3b0da98c534a5603faa9b984301c15edeb6042d7ba1171c4a1bfa08f8919e0",
      x"a5bc585e5c50e73c6761c4f3d59025d324beefdb59af4f1b7cebdbc9fce4eb8d",
      x"24e52e24e223abc807381902339d6d335e07b3bc5dc659470b5b31a662e18253",
      x"1b6567751d5bed14f050f6ff2f00f19c56add760ea367fde9caeabc5a75ca23f",
      x"88eb80e47126a5a8985fe2e6eca2df992dec34d342e2165fb3b66237f4ef2e38",
      x"b8c14fca1f51a873d7e082202330a3f825d95121789d22f2dd8c7bed9be9a160",
      x"4899a9eea4d39654d9fc989a03c5ed5c1de2a348c990fd103d25ac61caf0fb3f",
      x"1cf9b8e7f0cc45564c082067a81dc349f2f913b0f74fd05ee5b0f29abb90e8ae",
      x"eadc8924de1d1cd4473c47bccbfebae047f502030e31259293b53c4a9bf85908",
      x"68f0c77b345458b10731b6e38d786f17f7357ccd8a8726de6e163e3d3c5e383e",
      x"e2245a36fe52c55f292f4fa2c8bdbb3e40c2a5a5d32aa06add548f03e826a57b",
      x"901b249c8429c4732cf8308561b9097e32d98542701fe62d87884032ac5e1a20",
      x"ee751d625ac69f75fd0ab5cbd6ab3d182d04322f8d02c38885f2917e40626211",
      x"7d11489228fc852cd5e647d2d42270a1aad6c21f1f8690592a3427c2b1d203fb",
      x"57ff85a43eea4501171e6d1e54a06f38954b99dff364b7bea06a6715f8c47f1e",
      x"c19b65debfc5c5e95a908ac02f57ba531f12b6602a01833a00041bef720ccb8e",
      x"27989a327e803bab7c5c77dbd68c8674aae95ee50876decc1214ef853e729830",
      x"6111b283d83fdcf6059696b5e6d33f1e1cf5a39ca5928e26a3f1002f7098081f",
      x"aedf8dc08759b5bedd6e569554218894a170e151436d2b64bf258288bd7142ae",
      x"2a2bc6398943dee8f9773bb7b8d93a5821d8259215edd50d1dc4a2332eaba023",
      x"33d1173cdae510c3017d3d961583aa1b5c12042fd4527f7f5afd6533c165d551",
      x"8ac4f088ef62b4787f618ecb37b5a03758115567ceec24b3d543f50c7902cf4e",
      x"32a15312ced3d35fca836b0239398dab499c56af5a035c2abe14e9e81536c110",
      x"620a341fcfd7da7a077fef0c9b37892d1bb9e2b39755306786413e930bfdb668",
      x"a0942d24cdf971327a165fc8c30919614e97fda1aea1d8691513e83a11a864ec",
      x"5df1d58612cdc00bb97b717501ce3c5155a1b7e147cd575b959e7adaa340c236",
      x"d7117a680e7f8cc5017ceb8f6754b1a0739ff116ac9537f87b7a09a0db1cc1b0",
      x"824fdd3c21d107ed7dd4259b561ab17f036e33bfc350623d2a648f261e5b4d4f",
      x"9b17ffa6e82398bc0459f9d6e937e0f9d8304fdfea15dc5d795f9e0b4c6d5210",
      x"ea3bf4152a0405c6505db8a5f9691d35c9391d02e364b3bec250ea120e087ffc",
      x"6a9c06c78134b2dd04661cb5d0724b045a94033ab5edc6a9504b7696d0a6aee7",
      x"1b705452607596720084077647f751a18984b4b08b03bb9072be167184c73319",
      x"e9ce99c44f2fc564db99e71e75f88fd52eaca7b5a68b987eedacdb24e3206518",
      x"bc505af590de4d0c2d83feb02831c56e6583e2e111225384fa35270e10df5c44",
      x"9b625f93a66def25fcbb78b51270733ce58f8b2263838df4ed9d077625a98b85",
      x"c1b39eacba66981b0eed778ccd9671bef71b52a6dd114ae1fc0622736417f285",
      x"43c23e94804cd9a06ea4d341d1d4f7e7516e6896708bb2acedef27fba6f9d9ab",
      x"57f4d29ee7d64fbacfe218847a997c4202622b1e700405c9f1e6d2186a43d2d1",
      x"562785ae2f20b5baacaac3d57f7263ab5e97626dab4bdae901968dd5fc9f4ed7",
      x"03f9588541ccbbbd4276fb8f1ba5447f56afe2c7446bd2b2f494b9fe672ad3bc",
      x"b56fb7bc3a5e775b821d21e6f9b6bd7709f9d5a7a23e63bf78af412713c0dd12",
      x"a50a9c15dbf1ee8e2d1bbdf58c3f31a988bd94725ac5ca8896a413fe227bfbf6",
      x"184d51b3a1e180c43d2647a10113aa1ccbcf01f4622beb6aa6b56b1ea345dd06",
      x"7f84cf68a28aa1e6060996cc92b40bef1f51f49113cd902d7548006adc0138d2",
      x"eca21e2743964dcd6cc831ba67b3180b61eed41b908b6190e794dfa6a54e25a6",
      x"273e0acf307bb6521fdef9d59c3eec3e5e1b658b00a72d7c13791ed44fcf526d",
      x"f5ea8e242349f0bc92869627e0f05f83abc2a2cdf93a017c0b58f1ad805d4b07",
      x"f08e74054b380dc07a689d9b0f74bae4ebd3cef8b95e3b229546a2d23a855fc6",
      x"0c1e5efac16ac93fab82ca3fd6746a5f352b604e8eec88d2a3b7212fcf11e582",
      x"c607aaccbb6b664fc3a8fd47db29b927567f2cbba58f2d38a58bb1580f8ce696",
      x"49f4270605431a532836556416171edb67402c833463b0fc17ba9a6e14786f81",
      x"d610468d2386ff385b0b290fbe55ac8f8744669877de60118d965a2784bc421f",
      x"9685131c7aae5484709c9c31b5c2348cddf7f28152808e8c095cce82c801c642",
      x"c72a42ba2e33c3def895a5b4f19d30b353788a2b00411c97103e8faea8a16632",
      x"9ab00f957f27cb2aab6bacb31c19703711ddc55804fd12b6db26a3bdc2912a6e",
      x"0df3950d63e9746eb893eda5a8febb300d7026fad42bd3c7c004d3a3ec7a4959",
      x"d6897c6b965979bb18a89cd7728e1156192b44737db6341ce19f3a3b5c164350",
      x"4322023cbaeb33d517a0ff0cbc4c94c5c176b1a15505a374e710ff98900e0059",
      x"023ab8cbfb53370fd5f046fc93c1614884a96ca599ac92b51221c83b669229e4",
      x"39df7524c4c64c5c91ec0f2ba2be4ebda81631e933300280ae0f7bfb73ec1051",
      x"e69804058a96f4009981337e52cff0b7f5043e131910151eb04d0d0391711ee3",
      x"7176d842cad170db7157228e3285a203ccb2635a10feeb791a8b2cb8d2c3a35c",
      x"c76d47fbf5ede8e21f177d9fab87f2abed6a9cf3b91cbbc17f71d415f5c670df",
      x"9ab7cdbdc59e7326facce0c5e4800763f7cb484231912fd90402f47a2004f15d",
      x"595e542cf180afd78860847ada47a3c1201274a094c54a03d1ebf7ee5ba2d535",
      x"acf073b0a95ea95ef70bf830d0f36ee71a6de66beb26d5473a18a49641292863",
      x"1cbf83f4be0c6155b3db71172baaaae411cad34305f54e1c2dccca017c0112ea",
      x"ad295443849cee7daed0b42fb8ba8350e49b2dece9355e6c7a7f9eaeda8ad4dd",
      x"fcdbec77bc67c281d7e86287c5d73d942f6700e54f12edfd97dd1e515341625e",
      x"36012429c9d63091c83913d7b927675f3fb5927bff0581ee2533cd5776a48fbf",
      x"12f278cb15a6efbc453bd1479f2d2ccf21fabbb7f270344190244dc407483347",
      x"945fd8da0b275e29f581d5b55d3fa8df9f3639e6f6990b98cb75cdcbbc9f1234",
      x"aba2020c877e5114f000b8459e1d61312300984379cd880fe00d662b42f8cf1f",
      x"c1fcdef6d236914d35b70fc8ee8685768700ec7e5e2af364a40213a367c84a89",
      x"308717bc37afb816ac4d0ef44f8c7f8667a4cf713f7f17e9a96b37281efcf3b5",
      x"3cac3301f0f5edf51306f4f33d45199148aaae3712063fbefe8bedef820270a3",
      x"81132b7cbc06d17f787759cc03f9fa96d93fc4177d4c7817046f974065e8af46",
      x"a83065e0f90116eab1b2285c0861da526df755ecee2038cbcf3c4f87b82c86ce",
      x"932f92058d678e211df53e262db42642542a255cedd26c5a76702b4d9076c2cf",
      x"af1880c66a96f2f8c6f6206d59046c89d009d0ece95c7c6c5f4ed5969cd7f327",
      x"aea4116549f754a539312874b4cff06d23da85451512602e7006f2050d877141",
      x"4238d17ac5e5b66a1a1a2771f9a5bfa518460de81a4e761414ce2ebf6a844859",
      x"b53b6d6d733df33a6fa2739ba8be89d385ca02b0c030863ebc2c9331a060fcd2",
      x"ac17be69aec00563ab92b3f4c2032d371c21c6c8a4eae2fca162936ab670ab7d",
      x"3bfa118cad4259792b01b8c004ed3c2bf012746e76904ba55e3996bf6ca51f3e",
      x"8a51981267900bf72860ee66b747bdb7e1f0784246375e95cfdab9d9218f0371",
      x"9706cff1f628b8dae9260f18620e9fb30fb5245962299a258b7ddb26a278e497",
      x"cc5bd688e155890c3b635b815b62bed9788fc6fbb662961e41c01b5ccaeb0422",
      x"eff876b8b83abd07dea2b69fc6e331f5d7cc64c2b00227b573f839f432ed9b8e",
      x"dc4c951e9d8f3e361c6fa2f7eb2d6a3138bb3d73c41a12c2da484b5706db033b",
      x"1343731b0782d23678e39ab56f1bdac276f7489a1f8938f1ff82d5411f7b159c",
      x"ea970b831c8500113b7b07203a11903963999733afa2b76fdc4532f4ea6cdb5d",
      x"ecd241f03ce2ee3a74caad810eea17c26156ecce2c639d1efea52483f49dea04",
      x"19584ce91eef64d3c22d8a12172335d8ad1fd8e5e922519fb7b5deb2859a534c",
      x"a7603dc33ae4acf3bfddcfd4c94697b183f51dadd0211f2ad4a53f332aea29cd",
      x"05e1d7f1429c65394bf207a8ed9d8c301567e1059800dafb7714da28d127dae9",
      x"a03fce8a42179eaad79877156f4f20685c5dbd3b01708a96eda91e1e7ef9b62e",
      x"616e2a972e47e7e3e4443487e368caafcce394523fdf855d445c14ee43738c6b",
      x"c291e6e754069e73707cd1e1a9e03c988ff30ad0be7688df57d7fbdf96fd6b40",
      x"d4faaa3481d3f175f6de02ce78bdeb8402030ed63bcbf88cf51dfeadb3bcc66b",
      x"fcd4dd3e73a92516d68488d605204f5619ab226ca168f075dd0b23f26289ecc5",
      x"4f0aacb52478c91ba24d57ecd294ffd40aa6eb732dbd03ce758e058d9c8d5d77",
      x"f3caf980e3b9562519022365ece795e88bf42429915bedae75de6705a8e5e327",
      x"ab398557b177bbb7ac1b2918ffcd49d8041e0c75280d798b53202dc772225ad6",
      x"c80f9fccc84293c00a9e1bbecd9a66e7f467ecb59e803b3cf8d5a2cbfeddb0c8",
      x"3f317d47c488330993f5b3f83a8fa178b156cd3aac00d45a62c18c3cb796be4f",
      x"84abd459665d02c66934787fda0864620f9c122835b15b490820e6fd8ab6dc85",
      x"6907aa1440e5c6618017a044dba4c50fd546919148ea461ccfcb1dff8b9a92ea",
      x"e358cb266511735d8444c4d9a3948eecf8cf6062d912ac527db9a1fd3946164b",
      x"02fc4c898ec60f8c953b26074cfdd37693fe80eb953dc1659e58dbdaa0cb96aa",
      x"cc1fa696f6a50fc6bac1141bb40057d452fa03bcc51a5ff98bec5a9fe9069e4e",
      x"3fae5a197dcb7a3f13f93cdd6caaadce3627eced61ba117b987f7721d6f79594",
      x"55ad778dd688a6d83020f9699280d80e81e4babf77d09293c396a208262f8842",
      x"bbf7ef42258eae0e419110a1f316dcb52ac128eebe01a590ac8a4a120edb5eb9",
      x"feab4be009f1fb5cdd1556a84be303564ed0708c0a8b41524043fc6c39a32a8c",
      x"894115daa214a7321ce1ce45b31d0f20dc9fb0cfff0c93b9146b1e44bef70d67",
      x"486eaeda85f9a4b126c782109d4349855b51336530fd3b5fb6cb54bbdd87b849",
      x"9158c920c87daed0a2ed34c7ebaa45432d4a9f1365764c299df548ac2136a5ec",
      x"fdc473054c98efe7a998a0cd659e7e72d0f276861de27f0f077087f946641786",
      x"a62d6fa42f041be6ecc8b9bf4a8aa61853d36b3524299f9e5b4f4cdcc98988d1",
      x"c0cc9c1aca31a8f1c03a5a7b9b2254d8938fb52796493f7806dcd61673871368",
      x"6ea55d792d994582b4f42e396008b2618e66f3d05cb5450ced9d73e62daaa9f9",
      x"f966962a5637d0ababd24edbee368d1e32250e438a63d702f45a494d047c5965",
      x"0be84fe5eaca6980e41e34215eb1c9f6d9e9d09ca6533ad38b9afbaaf30c0fa4",
      x"e38b5fe5817bccf1bfcd750b0a8b1e849f64cbd119b4ffdcb5c3bae5fbdfc20b",
      x"2832f549813e6f920592eea6dd93e51a8f124cfab140aff936f565e239b2fdb0",
      x"ccbec269daf047f52130590ff60ab923f19ec683fd9d1eab49db682bbfff86e0",
      x"9fe57cd357a60a1cba61eee668f20de25a44ee7e0d168bd1f5380b0145cec3e7",
      x"06d8686fd3548b4e4e7f7c54d75ab2b8715515a5f0d08d89ed4aa855904330b9",
      x"f289eb16877946ad8d6dae205821047e66c0f31a4aeb899522c7561703cbdd2c",
      x"9c26b9850bb209af8512be0cc4fa319cbfa932e155879fd0c0074a1639ab6723",
      x"ea446c5a744a8471ab481e2334e843befeefecef485c561ac021521647cb5c4e",
      x"45e1c97a1cacda983fba8ca2c35c093eddf38db802766379cf6d73cbc532ca03",
      x"e1d2680db453aec385de70619f52b529c7460669f06f44abdc6a0fbce0001863",
      x"4c8291e871d0322cd396871c134f0b89c626a59264dc7d92414f19f2a75c5e4c",
      x"46dd0d54e5d98b9a3304f30318540ef12f242019bafcac9ec10da288be5af4dd",
      x"cf90f67fd76d3fc8c2883edb25495b8fb4e08aca07a4512457a5f310438ea7e4",
      x"858a1d9eed38f6b57d4c57a66df21138ca32fd9046d0a59323c114bde69792b0",
      x"3d0931bc41bd07d9c192d85b0ef3e02c8c2b3e7f455656fdf9a8ae53d947f533",
      x"46fa345382e53417b817e0df273626f8418a237c0cfa5921109c1928b699686a",
      x"ad6321d6c1c492b2d21870abda48d928c8b70fe64d45db00212d5bda4ee16dce",
      x"17a0482b803477db843597f063313355700bfcc24df3018f0c9ea0c9f3286cb8",
      x"c9811c6bdf06bfb6c61ef5dd814d85e0e092407f638f491da140f2d281570a0f",
      x"053e6e9ec46bbecbbff3f9211bfac5620955dc19170119bd194997a58c8c691b",
      x"31022a6447ae62de54f9a5811f751c197d38c8d3876db6f1db8910b01c1396b2",
      x"ef7afc9751fd9f082968b4363cd85d24188e434b731238263d47f9236f8d9d5d",
      x"bbdd3e3585296f8d69bdb3b099e03e6cfdbae4f25e3f39f87edfd2319dc19d7e",
      x"62ae036764a126e47c08c89fe59c6b55284fd235537ebcb4e331cabc7bfe7dd4",
      x"e4e194b824e90c0d89c6aecdd86da08ddab960f4458db7c19b382b4a7c55a8b0",
      x"b0e2c67fbaa68f00cd55d46d4e542736099d2ff22494674bc852465034f35ef0",
      x"8ca4df0c25dd261ba298285f107eda5c81ddbd88987282b020c00612cbb6e7ac",
      x"6781f760de43aa472f20f14d70a38058b5b9b4f12eacc2f164173730ac0efcea",
      x"5b23af68b77975023e35d2f7ab877b22f383796d1c8beff38677c3c3cdaa5814",
      x"637da3fcfd93639705b41ed72f8f642195e21098bbc68a5388c36bee402f1190",
      x"ea53d6714ecd7b01b9c3c5c934b64d7820d74da6576524e95b3fab08017eb391",
      x"f7b756519084d869f47c10b08cc27fffeb25671014d5c0a7e066a2b79c40f1f5",
      x"dcbc1f98e37597edc6cdb1c2feb61e547876b7cde1e430769c8b2dffdd66fec8",
      x"23e78e55dfd6dcecc8350888138281aab3d686597d5fe23469d8a6c851a2c04c",
      x"612305c4cccf25db52988ea1533e89bd1ca65d36de0a67da2520bd5073a5fd7d",
      x"c08b27ad8ce480de65387c90f07ea1769a3a3c3430821b26f324c1cf89449e48",
      x"ab95f549ec4292620724f5c6896eb70795c5aef141ebab4776fb89001ed170f6",
      x"024f30fcf169f5637a0428dff3e33b0ed65d15dfe66348e8c2379bb8b1faf338",
      x"f845c2a0f451df8e157a63277b7c95f235e0b5d238e23a415aa788b7be7fc619",
      x"0bbd2af2b523e79c1233673cab3b22f85ed522a0d77f489176fccfd245cef2af",
      x"1dd1e6c7cb73edabb3e5faf398bf2e678ee91dba2527ae5d89e7f84b78c4aa9b",
      x"4b636f606a8562c0c7bf190a868f55afe4640ceb126a0a571316c87d2ccafb4e",
      x"cb895f516c34a08f47758d87ea694d8a3c9a5f697c14c74703319ce2245a6154",
      x"70cea66241e0b19d8f0a98277e480e86942f31cd6d830d358a7d6114df3493ef",
      x"77f04516c450be06384e7a8c8ae125b0b74f303e99626f21fc70f3222a24e1b5",
      x"d5f5c0128531fc607ecd9fae42ab4cb28c9530aaac4596f2a4b1191fb467adbe",
      x"3b8ebf36f43ea163045b7c1112d8fefedb62928481165db56b66e996c5db1b90",
      x"795c8104464e0514729e62ef9c9aaa6ecd80a1e6678eb25f8ba55390f0c55b78",
      x"82b69072d3d9dd5c51d0fda5fa4834397ff6501caf2f53054b33cd0c2781b238",
      x"334c15b9604f2fc9a3640d83c4605b9ef858ec27f7c45fc259226f2dd54bb3a4",
      x"8c26508df3ed00a19fd41905e53821ad4ac3661d8a2f22eb9ca931b18f4a6b0a",
      x"a8461803919d6b0485b3d630af232c3ad764a200efbcadd3014a42beb0b3b137",
      x"211f2532f3c924e386c8f2b5d8d960346a8efe1b495c4615fedf0e844836170f",
      x"c930b8ca6f13345e951ec749d4ce5019197f56a829bca62d912537e6fd53afcc",
      x"b59d81df1521ba8d53e4542f08b51923e78ebf188e7e563f6dc234d7045c5916",
      x"9131f1a82826c70da011384ebf7826902a1e140a23e55ff766215eb82afa2dad",
      x"92adcd3b2eb6badbd51aa21e777a7edcbf42a8524d67445cf7ccdaca48238e24"
    ),
    (
      x"899301177b70c9f832e336e60dc6c7a38dd6065695475b76cdc64eeef1e4fff2",
      x"06a325b15b29ab7adb55c74e35dc093a1a43b88204277f5d6d04bf1588a84ab7",
      x"2761e25dd423b9ababe3e58d4adca49bf99cea4cb52fdf899aa5aa8796e29a7d",
      x"fc3577c78ab5a3a7755156ccfdc68720321e318abf79f45b8f73b15c0277c84c",
      x"485a2a831428d381cddf3d481bf10ecf42f85044f414c8d61beecbd023df5a60",
      x"b0c2f54c285ff2bc318278d1baaf46af176ba7e9a5b72465939d4d691fcd421f",
      x"a7c8b803dae1ce340349aa2f9c62819c9c00d3bbfa78ca8e11f894bf94d58993",
      x"4ca88b2da919e8f49c89d0e296b0a535f7f9a745b6f863a0779a365a438cbb08",
      x"093a1e9ee815077b1813b1e06802614b1ebf44cf9c61594e291e9fc5eba1f96c",
      x"75861282b5a9ca4feb1393e75817932ad59c63f17eca81c149ddafc4a982c998",
      x"5c3706b4c8e3e897573818d2f0d6227332ae9d24748ac694744c0c85b71cbf28",
      x"55002f6fdda12af82086cd78260b7ce6e9717bc62584af5d53140c3d188b6820",
      x"b7c0c6d0b1a3d39f7bd106e8986e4974d7958e09a332542c824e844b8f1530d3",
      x"ad012b00391eb4b7e80cfd0ed6c6af47d3755d9c8c87fd74eb52faad9330fcbd",
      x"262311dd9dab8c88a7f14c6d646ee98bd6deab70f80a7e0878231e51c6715c55",
      x"d42ac724fdd2e5e6dcb380fc40f1b6e34fc1d811d779b7ec026d2cdb4b95603d",
      x"f3cb8e82aa5c34989d4f3cb358faf9bdaf538b740cb8168d5c625c3698cde150",
      x"022c232d72c7a37a182ec8ffc1d65dfb556631ba2056d2a959da6ce3296ec9a5",
      x"b4e1aca982a226d275a333a2f233070873b2f341cfdeb557b95daaffc0ec8b4a",
      x"5842de97caae6b8f1dfc629b96a791ad0d52a0d9058a48a4227ff73a047cbaca",
      x"ec202b11edb204c1ae1eddb70a310848610c2c245b2b0ef093bc706b15a423bf",
      x"88f7c82a117c06e17d3d4ea30ab7824032082a01312c94e6198bbe77dc876cb1",
      x"d51e5e9c0268be56d1865ef697ca6501bb0e43e60f850b0b21a29fc3366d9c22",
      x"6fd5f36c98d00922bf3c605635380d8b16b90071a3b2a38189492e6cace95dc6",
      x"ac6e55466d0206a51607c2f313e64f11ba2575928345a9a2d10d78493ea6119f",
      x"abe38c407c6c05b25f2061fe82680a71ac29c4715ea3fb4f49467d706a9c803c",
      x"8a61e36e761d634463b1e58f61b02442daf0413b82a73a3c8d2cf796d360285e",
      x"9ff7f4a50f1a6a188e2ff20b6a18919f2ce257863565c7a77bb74cadede14be8",
      x"87be2ce309c9c02d1cbeb405898342d7fa6e8ebae6d059525e4e65c886449435",
      x"14211ab4687beb4ba95fa5c185028128609bedff9aa208497d4243660ba08bb5",
      x"37a5d4d05fe2d2f3b9c286bd9b12170e9754442f1b74ceb3e57e6c200956f50c",
      x"a044154ee2ea5ca8fc87c63346644281c7130c91e9affc4d62d02b961b28a647",
      x"58d67057178b496a70bb0c1c1f4d98ad09e3a998cbd845d9c2c10fd4d1652be0",
      x"01a808f92cb3b2ebd994a61380d87a34840ebaa5df05dcbc5803004172120399",
      x"fde590b338bb2cd6894ddbb53ee63547c802e407cc29ff5b276d8dd1e8b13abb",
      x"224e25f5c625f576a4613f30b5f24293002de17c6221144f32eee8871647f1a3",
      x"32698ee982ad44e5078a1e1ead3bd73e1efb1f0987de0bd192aa6049c2e545e3",
      x"492a51930e8be6f3c30586340c4658e62ed1bdd6274de7da98aeb4f56645746f",
      x"8436c5ff9c4818dc3045c2d1988783ee5dd13b34f06701f14243267c89590773",
      x"49479cbd8b58bfcb0d5efd56f825e818177adaa88a6fad814d99420fe8fc4141",
      x"5c100e281d3620334d7bc1efc08aaada9f0675207f9204317606c7936057375f",
      x"8962565862687dfaa7b4b81705274e36e2ebd65cff45b6f0a4b77ec0ee34d447",
      x"911da380b549f2a50913fcbea1994c75cd83ca6d76016545b63d6d282f48c64a",
      x"aa8e60d0fb091346ac94de1d0ee3f5ab4d7a4a29e86e756dc5af32a0701e8c00",
      x"b4c3027e16009d8dda7b20db12364990843dfc2c90067fc68e75ae353c70c785",
      x"8fa387b2a6b39284fc1ffc8a7c611bf5f732a3bc22bf83a24dca1821b1141019",
      x"1b09c68ae414690c56b3f21f22cdc4010c3c0ac6df39267ea403001c07e9c798",
      x"971ec18be5dadf4170fcedc0566288ecdfede6e3c3ff7200c2eeccd8f848abdd",
      x"5d12b877d3128761672e80c94d20420e5eb10e9ebaa42a07050469beaa11404e",
      x"91e1b92f12109fed9417bdfa9904673827d088a8361e34e9d2c216f4e54004a9",
      x"881e7d5ad74467f9b7400d99f37f0a8e73cdd68bc0d6b9d08a673bf01fc9f9d4",
      x"3ca0583b50ae18fdd0efb8c732d1a2c9f7c34f8f31aaf69ddb96fa0f2c91c7ed",
      x"fef2c10cce743d4592d93941f85ce25116e618cf45633c1f6a742ce577c3bb05",
      x"dcaf5df78c754bd2f16415bed739067b15df7558c8b436af37f2e38c16a2d3c2",
      x"ecd3850f92239d84f272888ad4063ab30174882a8ec78c7c0b5feb20ea8c6cb1",
      x"89304e7566638534bfa4a7a977aec362495d7de7e57b568f1114c38f40930fcc",
      x"343ca3f79ed3b7c1cf2f5f391667afef5a9c19529a5860ac66e996166fd731ce",
      x"c3402aa460c9215d71db2c7d005ebf54f7fff4ee3bb20d6ecb26ffd7f9762b93",
      x"e3f2d2d2004e0cd897aef0db291ae98043586fe5efd3391fa53af242311c8ef9",
      x"cdd1f8b1f6a9ba6430bfd6747e6800058fca772973beeb069a4aee99c5207f26",
      x"2005d1600f843bded050dda421488b8f80cd610a2bf6163c88bad84f89a14a74",
      x"08fc999fbd250415fbebd167cf0ec64849bbdcbd3d5e6c9c0638f2713a14836f",
      x"061ad659aa1e03eec470a53de11195e0de742542b6895cbcef1e81b348c36d46",
      x"bc85736d5c591d900673beae65b386d9042c67580b245f9cffe1b1ce35118df5",
      x"43ae6c2a96101be42d7f6cef198963dd21b11b30ba3167f4ddf5257d412d7fdf",
      x"db7e1081afb485113ea09ab6236a0a0f983f4a1f96b6d6ae00f88ad792213622",
      x"1e93b497db5d57327b76eed8423ea4da4e77f6648f99b0612b1e7561cee94e24",
      x"8b3523263dbdec1fae95856fb119e6cf5a4b21a5cad942c2e0b71c1ae2c49210",
      x"663ffaf4bf1039b898dfe5e4a102be546bb8a861fdaa56008fbc6ad396fd12f5",
      x"e995e1a9800f7c0c4cf44d25720b7af12e51d3367d8363daab7fb6cbdfd2e16c",
      x"2c25f1344f57ce0e7415946d20d7191809b87220763bc9592ab96955f0461cdf",
      x"bfe74d6189672f101751a855ac1d12f080606c00f9c194b99dfe09c2825660eb",
      x"44682dbf52fec5b7a3898719922bdbd788293dd3e738be939490254117297410",
      x"3d01f4aa9a860deaa8c5cf25b1f12add0eaebe5ae85cf4861fe0a4dc2f12ee27",
      x"5ff644a0ba1d4bc4c42f3e9d12739e5c197326be6b4498505218d95ef576cc93",
      x"fd4f0ae363cdb82eaa320d5237a8cbdc366d557a1c257c078f4cf55d81cbe992",
      x"0a1bdab1609530f993a8e06d04a971343badad839974c01f9b35559bfae11a96",
      x"d9878b2541c720e030e675724f1e24e2bdbaa2a7dab0a27f2e33d28aab01b371",
      x"51215ec45062998cbca6cbcc31071c39b9ca287aa7fa2ce7e1bbc0df69e6ad38",
      x"52af3c2ab5938aedce5b4f0e80b804e01c2450707d1558c9f5dd67276092b146",
      x"26764f16aaa146e52463ee779738fa32ff04ff9f864e06acec35c82443a08648",
      x"55a8ea5c0a6fd32a9b769e3eb6b34b02197e459f44f52ef9790be285a483d58c",
      x"1184db2e9e3ca372b6133aac76097fa2a9f00dced626897d24c2f22ca130dd88",
      x"824655bf27150220b6dbd28721a3256c25c0234820a09a03b01c81f603744009",
      x"db6abd4337266c0b72ad5641886579c885194e4cd9e77555b567c1872c637bf9",
      x"a5a41469996bd9e2ee33256e55087941541ace1587b73cbf29d4dcc90be29f7d",
      x"87410b751a74eecc880258ca95490810422d616c19d8f16d6eb10e7721439c84",
      x"09c200d10b66f5512908c9f65a844a32d23ce4f2ac7df12f5550c1fd135c0ea3",
      x"ed9ae8b229e92ee2971e0548db4e5fbce15030abba80da2790d4ab3362c3f9f9",
      x"e122c78d7c8d38465819db98693d77a205fea386c6e9c49863e0a3ccfd6ee909",
      x"68e4dce13925e97d4daece0b8c3d8dc427ee10f82149717953a12ab4326baef0",
      x"4c6196d59954ff448bb0a6a1abb7ba9c74177d41f298f16983c9404caad249d3",
      x"e1d22d26516818a463b40e3f83953567c289b39bcaef6acb56ae46c6ccc3b606",
      x"4d5bb3988df1b26d6c2ba7a4884a796a2c588dc5e84c17979f449d6d3a682847",
      x"bf5b4c8aa06896ba80f682f4b49f78aee65485b5488a5ed4be721e8a1b0e65de",
      x"8eaed96cedebf8cf9ae671e8c71b3124e792eb04bad0bbe8e6ce506665b88d62",
      x"11fd438bfb59fa2f5c89931072a28f7a72ed881299a7fae42e8130961dff5687",
      x"348de59836b2c95a263b51a905b19ab6a7761f4c7730d069ef3eec0d4d785286",
      x"236f65f001f3402ed7bdf70a015d45ab5e4ef5a44de9ed88f15431c3a527b9ca",
      x"dd7a3761276dbc8be5b469a77a0fbb22daf6edc00bed339e367ee93d7feaad03",
      x"8aa12a26d1dde252af8fda09aad0a1d122a5a0977dd13de6d4d67fd48f8fd860",
      x"f72ff684ac45a71f65a3fa670af88270d4397da890eb77eca4c38c401d62e33c",
      x"55553e9cee9e75806b4d6067d994fd1ad5f6e4f4d703af5eb48c268946b490de",
      x"9b8d7a4b489defac6ce0fef13643c3960c47faeafa4f395692c1e85bd005cd8f",
      x"cbae91d9aa6a92b54e8a6702cc8642438b6fd2e32160dbdec9b6198febf4d650",
      x"8d3f6c63092e6a3b56c08304e926b0aedbffb1cce5d14d3c4e21317f97d76d0e",
      x"ea2cca71a7132bd4594d856c0026d11f48059dae44fb2407ac3abc530f9de281",
      x"9b2479de5a8bc698481e011b76409404b804c78fa5ff5d813d2d0f35ddff1027",
      x"b33b2801d738efb7f9e65015a84d6d2a2ef35f2c593903bc1b05f7d8a4eb1f47",
      x"86b0debd63557830e5caa4ba0943929871fe8e535c6b72b6bf33c3f8124619b2",
      x"f1a3de299a618435c5b8d2568f17af8378ab11d17027f1aa80c2eeeb33929afd",
      x"755a56e833f0a3ac1a24e46741a463e98ab90aa5906cdf702f75a3cb29dbc4dd",
      x"a1a8e71c99b199561d8dee62cfb83767ca3ca023688235d3c7f69591da7a3061",
      x"6e0f4a5ece8e12829f3adc5118e9016309899b99b3184259c52a90e4dec29bae",
      x"e304baaf9fb2700f10a36169ee6a72eab561cf1d1d9ed5dd414ecb3755e57e7b",
      x"3c422640ca0ef466a48bb1e3bbf27604bcabaf779a068d753da8085a933e37e3",
      x"a817b904f52cf6aa576e9be18f16a42947c23265d9e5b4ece3a76d910d2eaffa",
      x"f582e63ec9cd8d5803612112268614529af8073c76923c69c0347de468de27a8",
      x"564218bec9e51034b4b1107ff8d12ea57c4d772512fede23fd70db13d408dbdf",
      x"0dc67d1742c074668efd7278e47b1b579ef3c6f0670f0e209b075eaa14ccbde5",
      x"fbef48dee557f1129135b94d0f6fc465c92e5b9babe3f65e29ff69d0256c7475",
      x"ceea76caf9b63a8a00c0d619aa66c391d022a787bce2b824a8b4eff060ad1fa0",
      x"e7d3b8467db33230fe4d0ba6bd65269f482eb943edbd279e8baf90084966c5dc",
      x"c1b4b2995aba60a70d862c6b07ef9e73639471d3879ee6de59567fefdcf15f17",
      x"281e6537d35e4ca0155fa1f4d9457c31724f8a8e887c1d510ea2ed0ed70d6045",
      x"70d719f176be9e3c78d326146d04d7198d1ab453c9fcb301413c548f01e5f0a4",
      x"80245e716f4720e86a643f4f42165b1ae32e88a29900b2bc5335c590e48ff151",
      x"094661332b2031d0fb9fd67971fda16c5d1b8e9d65e63c7efc12fb910633e127",
      x"eea79aa318323d837e02b5fe98e0801e89ef09a301513e52c335aa6ffb936e22",
      x"43f7489161213fd96cdfe437232423e5ecf9d1b1c87c5c698a9527d7d25eef49",
      x"0eb7990d1c2809f95d8c3d92f1da0aaac30e2e12e78430a837590029deaf6cf5",
      x"1938c6c2985ad94310f6b6bb7511466a383c6c204147b0aad5cad9bb7b87c59f",
      x"2e39960a9549979e86d7895231d754797176eab7e4172e5816be570c5ff73b3c",
      x"13034fac7584626221a003e92e2f5ece8707a5781d0decdd6a355473b965c621",
      x"55955550b491f08797c9f17fc8d73c55fbf0b237e459a584bccd637a720118b0",
      x"0eda68386e599013fd0513136ad5379bbdcf94cd85cf775974b49c503f68e3eb",
      x"d29f05e7147085a50d6b17bb93e6da84373f36acbdb1a1080363ba0d24219ff0",
      x"e5feac794701100c9c1cd3b4a1823eded8723c8b6737f7cf76657af021a1c5f7",
      x"6cc43c6fdf327a36bb80447ad2a76b5367077103439a762c5f9e5ea4de2e43b8",
      x"bfa9c11266dc78ec5416b8dd4156d32d3e4b904b4f2855915f250c8dee7c271a",
      x"9e3d137b089cfe45e21f79e2506e1cc458d45d48cd2a7f94f9cacae064ebd0b5",
      x"12bd08c694640abd38a75ab4f8216a7acd42cdf712b567edb0bd61cd71c51f05",
      x"d9b7ecd5b14d442b25b8ff1b10c4ce44dbb80e9e9e6737ccfe567806c30f3a97",
      x"ae6c89cf4e089677482708669505faf7c90cbaee4a9afb9bbc98a9d59f9c6c20",
      x"4fcf202e13a96b0af3150a53cbef20d1be1e428f9b6017856e64ad40ba50295c",
      x"ee5f989ec922eb3ce26dee0633a7c719648371321bcf38d7a821b82754c9c0c7",
      x"2fd24a7647a8a456282ab8e3328df885c7897611401c9a2c2e0cc1697da73bf8",
      x"2ad9da9ca136ba79bea3d622090f56a11cf5db0e5e07fc2f4d9bb90ccc1b44af",
      x"f8818c70d6b4ae40191bae9ba3d519282bb7738c40dddf5da480d541426d6082",
      x"7e916b8f9d254f0c981103909fb032018b9e494c4418e74b3f4b49975c9f23f6",
      x"4cadb52014d43f1c400145fff5cafd4e6b6066862480ededfca464a85cd98640",
      x"8e868c0f1806fecabf1f617f0a6ad422d506d06760c2860b711ae2b6f8098de2",
      x"fc0ed723fb1ac2ad486e327e9b9b0ea4bc78dcd82e7106f26a335fb7a7fae598",
      x"b170a39d40b01566930a8c9f2fb7b1475002b8b9418ea7adb6d4dfb8fea517aa",
      x"f3dba23888ebb2019fe93e99dba6017c37327620aa3d80b995522844e8138769",
      x"cfe302095194544b22a4ba7abf7beff31474c0041f356d115e02e90077fd1b08",
      x"006b8416b1bbae745ea30961626138715f70bcfba87e17f988c4bef867b5049d",
      x"541f949545ff6ccd80dc44f77bee7b25a31db59630b706356f281dd0685601d5",
      x"b8bb500514bed987b8f50c21b87746a225ae98bc57a51e7c963b029dac54f05e",
      x"e57bef5070261e38f4ab1857bdf88a6c0ca1f75d62b86dad36fc53cb8f7895d1",
      x"2b1ec356f4cb48c24aa11ac939abc99114b8a7942d7c6962b3ff64dccb396610",
      x"a63bc7495d43efac676bd3dbfd89dd292ca1db63e20c377d7066f841e1a2da7a",
      x"716d220b0947b47b86b970656156ba5c4b07ca198aa7fbc58481c68df4b78714",
      x"fee36ce20568fde5956ac04420775ff4d7be033a1e2a385d5cd34bad826ceeca",
      x"efd0aa290c45c4ad071d790545c3c6bf6a194aec226d691d0ff4c51a47850d07",
      x"040a0284accac598c14c52383e6d73fb4234b26d3df11cd9e3d0051ec4b4b12c",
      x"4ca05de26b5d47e3d6783389649b9085b616604e331d312ec27985e1b742363c",
      x"f0c26644e8092fe4af3f52af369fca03f00062f8a45bf62f71f7252d617b0a3b",
      x"69dcfd4081c027f74d59d8ab1c79bdd71f3345ea0d6ea91a2c551de52666d5b3",
      x"b5a8acb801ff0e57dae30e647d3332d286042701e975982044906a63583138b7",
      x"9af1f7261e9af6ed761d55289e871f87f3656f229c02a652aa594a2df2b16d07",
      x"54927d6e35d3609c2f92c3eae0e434abc4827011b7033002a9a62a996c0d65dd",
      x"b4f2f2adda55c7ffeaf8c6bb9f87ca0fb3afe7720b2ef87813aaafaa02c31f55",
      x"c9031a37599de2445f2e0d9515ea6e7ace0b727f0a0fe28478410819c6a74a66",
      x"213418cb3cb04784662146caa1838dac108d2379a17147f9e9b9c30552281876",
      x"41922f94caf2643819a7d0df59d32648a9d9cb2281f4367dc3793e5550dc30a8",
      x"f6bd82868cc6615eb3afe1a53938cadb4a62d6f93e761b8d30ecf309dcb53dcb",
      x"711afcebddf38385b86b62e85c8d7255537c994862654f77e72fb6514198e05d",
      x"4d678d2f57d107fcb2d25dbc92564f04d64c6adbd16725255cc00d82f0339f99",
      x"3d5bf83d21152637c4d3a3f0569d785eefd06081d42ec584e8b282d83e62ef7f",
      x"cf3f476a9044606d6d999983d02abeec35c5f29b20a7af9ce99bea9d9f76b675",
      x"cae4de924bdbd81ece8156f898c70a9962d3bc289a689c308d86306ce27797b6",
      x"f3ffd3942d361762293eee4b0593ff0e6eec19966524eff52d9442f5fa3452ec",
      x"b388e68bc0b2a0aa76c6b583d7556c9a794707e60c6b45171877fcbcd95d687e",
      x"4c9a39ba42e455099088ebabf423617fef2b61742fc21d43861463c6de2ce968",
      x"4aed41257ccc819dd3fc88228fd2a31a5e86affb02e82d1cef2c9dd4a6ebdfb3",
      x"5989eeb8567ee4d238100ef40c481dcc0989087f28b9a1f494db7146a9122ef6",
      x"eb67e365164eac22099f5adbe50b94cb2734bcde146a8b3eb013bcea52d9bad1",
      x"23660fd859cd0dbd58acdf652d2ae0e3815a008f93ecc6a17fb9e810fb29c7a1",
      x"e6b6bc61dd14f9c8caa816b64bd6c2465b1ea35e71f790988ca11530f788d621",
      x"f09720f7980d3c935aadf7aa2ec29be13b4f72494ba273fc359b6ca6bcd5cf7c",
      x"751adc4ed36bd84ae04c1700e6403c85e1fa8a1062c528d3c146753fd7f59517",
      x"dcf1b09b7b14f02a8bd1bb84558ca2f79fad175dfa4c6fca2f00a4ef10379d65",
      x"525423d898f84becdde6e22ff52ded69840fedbfc7551c14b74c5bdf32cabdd2",
      x"6aba99b888d7a013b984e9569f30f37bf7ee6eec76c53e7c0553babae68c7bca",
      x"a0e160b1e31d8d2d920efbc79bc057b325a2c4cc09a1d3e4acdfba282cadc6eb",
      x"21915846edb7c2b6e858a34fa0c0f6e7742fe0d4faf9a757441a95294d1b535f",
      x"ade9b7a52ca6dbb845031d631d288ac756ea6d591e8e296e3d60abfede560f03",
      x"cbbdb04f24c11eab9304204aeac8c70480464ea7075120cefa1f2c3c0cbdcfcc",
      x"6c1bf89589fcde62cec281f234281e67bb1094d023cc35eb9b4fb84822e7fafd",
      x"6622280e19878f5df85a925141e56c009cf0d2646b2600af62cf85458e6cda0f",
      x"3c76077014aaf49115de2b75b74045474fb8386bff82da62893493d270c3cbe8",
      x"5d38d865d21254ee0086677cdcc45ca14fd0bd7dbbcb5ec8538b350390e268fa",
      x"c0afaf51de865fca827bf82d2e125743d9f2fa24193c21d8c6cf7cef72fb4b25",
      x"3e434c5fe71d9c05f479a0f4e418e396a290f64d780674707c5d46f5438c5caf",
      x"8499fc47543cde52a785da01a54c40d54c12f011e698ca192a14b9cb290c677b",
      x"95759b322d035140f42f9377abc0699e7ad8d9bbb52c1cfb709f72d3e8a05cfb",
      x"fad8eb8bee70f7d2b3b1f94ca4a4a40dc610bc89ddecb96b7ced31dbe472360e",
      x"0c8cdfd55fd188a8e3a169975a7518007a731c77694f70ba89dd1a781840bb11",
      x"19b35e2496023f39589cf01480656354ce46556cb7ac9c0c8e29f49f29674a04",
      x"70d840f09578c1ded4ded80495f69c0530154106b37cd5e9f3fe0c52085cc058",
      x"ad376ce260120c5663705569afead630f1fb835ef89bc81be4060e2be524cb91",
      x"a4001b324fd63f232adf509b2c58a550eb711d2d6d6d4279a93e1ef6a32a9ee3",
      x"943301ac4d2d64c2543df75cad4fdde7af4f9efcd0f9c7e44bcb2416273bce5f",
      x"8ddd01e6606eb69ad3d23fda3bdc00d22a4845e2af8c6429074a21f5b62437c6",
      x"478d4b99b98332d0694ccf05ba719f6d076cc9501dd7ae44f0d594a56350b85a",
      x"3a5ec179a245a9bc0b6c7b45021ff8d4d8a5683b3832a4c88440fa468a109578",
      x"3c13791ee44285b9e6f78a01337f7e2e2739f747486c08b64ce92531e4c52ef8",
      x"f1effcdfb3196df215e89865f86d79ea1811713ee6f3894351b0f7ac86d8cf14",
      x"0e3900fa57e298cc3d11ede533f52f516e532ee5f776dd29ddb6ba0c886a9cbc",
      x"ab290ba95454fc49d9a0b86f5be566f9c74c5b801f68d94999885978da9a9e96",
      x"fbc84e1b9c2f371cbf5e964fb4d18491974c7a1e2ff41bf180355f0fae6cb542",
      x"80f665cb1fb0145f0c85b5e8bf0862d26db5676a5b2589704f5e08a1c2457802",
      x"1fa01e8e75432d151d2c3e6e8e3fd77f65bd9aa8b6e9502e9d1c99bc9847c616",
      x"5845e8bfe4771f9c10e4e5c082b3150af70833e595548f300b2e9dfd7f81b03e",
      x"bea8dc4fc67c7c2609cd233fbcd9e91f7e96acefa8a8aef7c1755972cc36a77b",
      x"c8a284e8ee40b33c2707207fb738926992e9f3e4b9c4c375a461f019d06916e1",
      x"54756cba437e589426ec0cc29652f12afcc4acb93265ebea8ea32216d359da6c",
      x"891aad9d6f8b60f1b9bf8bb085c46f67df0159ae24819ee0d6db01135fc40f6d",
      x"648cc6f510ae80d06f95e42e80d927e98288eded4f6f7e38da66e994951754b3",
      x"463399225ca0a7310c671174c53b1c1d2dda8ec364fc43b53a9d44d25605a015",
      x"5cee0ec706ad36a5983110fcfd29bf43d506b78cee52044e9fe11e94cd847417",
      x"4572cb0ec654428939a6d9682d19264b7b3dd95ed9fcb70ba3da68e0d84221d4",
      x"d076d735fa27cc02c123927faf1264e0aeef020de98a7c90412acefc1340f87a",
      x"296ffb647c397bb82b95039eb06c031d6298b52128bba11c67e2b9b0aa69f322",
      x"58f85d41db2fcd85763938d3b380ae3c89b7ee1f3d353fb7662ca45c8686e8eb",
      x"9a6d67177be7991123b95f66e7eebfd170adc51eaea342bd6f0a088be79b5bff",
      x"a7a69e8ae207b594ea04ed5ac99c0b76218f7c7a8b73e1307569dc23d7dc5b4c",
      x"4d14f77aa08b8fa81865c61d67a78094c5f7278cc5491eac12d1e41062b23c8e",
      x"9630d383b70b2fe840614e4a2f0e08c7ad4cb8c660cf5ed8882923d691d40835",
      x"39bd3dedb72721353b8bd6e8281da4f1a55aa8783f0ae9cb94d672781cc012d1",
      x"5c43fe90b521ac7f2efa286d5a0bcd2aa17bea1a34b5fe88844b901ae928f802",
      x"9405058cbe60ea89a68dee68a3ecc2d29b13ba324d21f50aa18c87a0e82e6dc9",
      x"c406d22aef21e248d070f329bf67066746aa89b5fa83e0a619bb787847431b90",
      x"2ecde76aebe80437a7d72775799f07e31b51cbbf8c9abf9148c1f530e3fa0531",
      x"b9d6bf093cca265661e1a4d7ca3595010558da76e11c4dfa8fab6ce1c44d6078",
      x"d443a2a85b2bcf0a5ce791658d3ad44e4a29e4d1a221ff17bb2cfe2ee663e879",
      x"6883acc548650bcc35e66a8a82655fba197644233fa221a6b9cdb8c613b539d1",
      x"0938b21b3b9ba41aa22322665e8f7739fad70e860b0ff31e4e3aa6fc3d264ae7",
      x"2870e99220e52e763255fcbae2a389f4bcb3fa2fc74bcf1c4bc14591714eb3ad",
      x"ebe5482976a8df7bb7e792230fda1ce23ba5eba78142b89afe870ce7ad57c826",
      x"b19c3ef60df5dbd8676c2f7700395d86c730744338e7b4cf2d0af62f32d7e6e0",
      x"62ca07d113f1006407186901e5cddfcc03c18a73ff717eee7c730dde482616d2",
      x"0c17c85b263f5b34614ec2531e45e0eb5fee9425d4ab82d7cdaf17786c22c2c7",
      x"30cfe7e3d969dc82f8410e3a649efaedcf93cbee42b6163ef0287275501a77fd",
      x"5da249a28a6be0e70719aafab3b39ddb79abf119c4456d6add1524aa551d1c60"
    ),
    (
      x"d9562217d970ad401fcdecc4541a33f1c8727f3abe2d69eba4f3666bd617df54",
      x"1514e0308cb14850e724b261b9858515539f789e542294791a750f4aac718cc3",
      x"fb0d79f96e0097081c5671f19f64a3f395dd4711061721866cd03eda224560e5",
      x"e5b50b165ab2d43bf2dc560e26614f057d2517269349f2721c7fc81db0bbef0f",
      x"c153f35748a0de47393a6ecd339874ea72c35b5b18eb335a34fe58f1b1cc8c9b",
      x"9de559d24c26eb1e3da0bc7a5dc16d8eb80d102fcd6220d20403cb7ff3c79591",
      x"f5c2f0bcb84ae632bf80a86ed9597c2e5afc02b8d0ff8daf4d42c6808ab1a59d",
      x"a0aad1e92ee201810b8f160a7cca25bc8d39808fa9b30e9f58dfc0e77ad914e6",
      x"e809c27ef80a7f27864377cc778ff47cb23b9de33edf296e186e49ef3af15103",
      x"4c95bff8fc85d33245176b53562899ecfd5d91e163322ed41c1ed885afa7fbe1",
      x"2ada93116d32045b8cc2d07b16e7af7a3113ceeabb2b6b7bae91aacfa3f0f6ff",
      x"ef3b4bf06f5233b8524089e9fb5c4e3f782de475b94a9bd14171835bfb8aed36",
      x"48581b2ee5eb0a9446124244b3a4a97d57aaffb07a5563f0f4dc8ba850d2f301",
      x"6e6aefd6a1c3d057e53bf0aa166aced923858d0d35b995bf1266ccf2019d2adb",
      x"b6007f89084ababedb855b3780f1ed8235e522072f9b5be2be83940fc341c866",
      x"cc80aa8152fddd2ceeb8c455fcae02daf66ecf10a2304742557dd176df13ea4f",
      x"efa5f121e46ac9f470735b3719bb8cb57b4e41c68e0e504b2e34cccc05cf3ca0",
      x"2ef6546ebd671ac200e47990af4070b0ab5b48aa33b1a2e41115e5affd90aa84",
      x"63df0b579b7b31e5d2d3c667b3af1f9fa16dd79c66729e04cb9c893c54e1aef1",
      x"80139a1fe2386451ecbc02816971df1bee5479f34dc173e1ed903e5ecc12b97b",
      x"8d7cd5bfeba0874d28e9d46230d0fdbb473e8fa9b251d3b248d57ec7da4954bd",
      x"852d936f11efe184e0b7ba37202ad9a39c5ec914d905ecfe5fe87f8973dc906d",
      x"bad1dacabd35b78e572641000fc3c7a52d1a4b50959fb1e327445aab6205a936",
      x"616f1c1ca84a9a6d3c636526dad5a23c8837ac845851c2fad0f54109b817110c",
      x"68af81ef73afaa4d1aa2ab68db12f3edc7da2ef113a6a6ca63b5966f08e77a66",
      x"98a7f5147515ea3d4f0f74b8b2c4d1267dcbbbf77b63b9b6b0f2cd2edd53ba29",
      x"3c5c7a2a23eaa6bab18a969a83acba08faaf65a33ce3916b88951e3bf0ba60b0",
      x"af8e94729c56ef1b7e6848b918fc74ae0966a6eccc65a1aee936aed849d0edfe",
      x"75cc7c86dcea7b4ba6af8da1b37690bb570364faef9a0ad53df20aa4f3974bca",
      x"9cf1f40ceb6be8cba14de3a7d994abb6c9e7923d6a12839778d4177902a49c79",
      x"a28947c5ab5826f10f7bf50a5a8615b2da22dee7db44deae943ccef7f39f01df",
      x"6ca7966fbdd04cad21a4d8a17ab1acd4043a66b29d93a59d057fc0a83743e9ee",
      x"01b9138981ea895037df976eb94a9c4b109458f594786e5ff951bfd81927ff3e",
      x"f20075c094c959f2b595b0316dd88291a933317c8b755c1dc94d43b96dc75282",
      x"d277ed574bfee61e45c6e4ac6e161d4095fc3c26330d92ddfe1da2c215b462fc",
      x"840d9557e2240936020c53e3968cd7f7aaffeeaa24c563af2f5f8989f0bee668",
      x"925a4fd5fa2b9e882b1d14edf14042bfa595bbcf021397094bfa68c8b101ce73",
      x"67158aa689ba61bb8f64df006b306e54997132dbe70563d25fff9c0dc6cfd4b1",
      x"6ee3c2f50487b0f93fce7a7dce5615b78910775c89f2664809e0ac392e752a93",
      x"3279fe0810afa9353d2afebaa959826f2f0dcb17b637ece6104d4ce1c0957df6",
      x"ec0b00afe79c5ea4cb7f8a463d05e00c736106731978a396ea6a7ec86a9166f2",
      x"c469f39fb7cc13b1dcb4e3e239ba92859b601deec88a3be186207d863dd8e85f",
      x"7dd716ac29b4330c826b56510f4a4e982e3204ddbc0f94aa322630e808c8be4a",
      x"d3b740615d7f46fb84b283c57989e29a703cb83b7df4516bfdbc71d395fd7b50",
      x"90e59531c5a07678e8aad461e060318e96ac208b54358b43c736699989d5834e",
      x"a0a30899a7572f055d9cfb515cf394b42abbb0414c1889f3433ebef3fe0a88c8",
      x"b983eca1b4527d6b52c23df0b48dbcfebd73aa5f07901e2108571e2bfe37f40e",
      x"9a97b7a0a9742e8ca2f699de83f6d8561872261020a439cf2229e5bba0f84dcc",
      x"79de6f2b702241d2f7fe2430764d9b5bedf7793d74491e82d2ab62b274b3b62c",
      x"114efdb76c50fef07d82da61126626da42f05a0cb455f96b674fcb21d0b0899d",
      x"6741d6a41c3238663bac51202fd83e135b7d80eb2fe48c06f1c8ef3df74cd4e3",
      x"c336aa35ae948da455c79ed7583abc3680e9127f8dfd50870acdd7ad5631fd8e",
      x"e28f9cfa1d44a56e69dfcc2c8a56408726dd27e72753db51414ec6d7e6d1d136",
      x"bacf1ddd0e6a1cdedc9cadfbf4f02b1ece0cd73e6e2d9388078015afc5cf6a78",
      x"57636645902dc245fcd0f6fd3cf3f0992cd9302a5955eb7e8011b87c53c11473",
      x"a62669f53c32b23801cd4d205ee5f37a48a74981c6f1118f69a5eefd5f507024",
      x"e0ae9bb5ef863af06dfa5c02985d600d77dc44696691bc8df6b94727487883e3",
      x"fc3539b147cee5b40b6843254959106275458bfbbd6b7b70fd2da73bcf0e6354",
      x"0398ab9823758499450b761c4ed58152351ec02d68bc94bb9843482f3b03620f",
      x"8c54e9ece651b4f18ff850ed270f47b4238cf8693e0232ae1ef182bbf53138b1",
      x"6399da01150a6762cd446e4fc27b77391dca95d4378ee60b2bea5d2ba5314b3b",
      x"fd0e882bb07a902e26cb4070ab3a95d84fad2b6d8dbfba803f33f909655028b0",
      x"c5c395638c3ddc10832aaee729b1c777c9847864173a829305ffe1cd571fe29f",
      x"5f5335649fb3c01eeb060ddb981e67381f27dcbba2f4b5cb76a6aab6030b7ee2",
      x"18c4b875867b333e1af89ff5490da9af5dd1a203981d229b469b0fbe7ebddfa9",
      x"bbe87a9559ae008d88afb3b3c2f577a92b879725b6f49e7b563f909b77f5c616",
      x"42b3d22f40da4e1e370ca98177365131709440e9f1287562cc68621e85608bb4",
      x"5e7bd9f59433244535496d7ed63754826bead4bc1b3bbac38514f1b9419e3a4d",
      x"74be11227cbd65714a7419e09e2e69ffca1ea1455a65efea3cb81c71acb02146",
      x"77e94338ff23b5e108526ebae943c5bb4bdc98857e68e42ded825ccfd65b0a11",
      x"c844cbe4002991baddcc7d35dd68dd5017830c6c7f61dec3c0b66926997683c4",
      x"f1927e76ab423dec1ff5f280780fbfb9c22366dc0a4e54a5302b66095eff42e0",
      x"9e66ea33a79786fedc73abc6508359d0cd2457876cadd214bb723bcc075eec90",
      x"a6fa7ae21497bf2864351f3811b7965706abf05561dcabe47ebd10793432de53",
      x"53d77ced31547e16ea538bc02dc464779d78d57633b38b7fc016f00af3951b3e",
      x"54f49189a70a8c87fb2c9f158d20f31d1d4fdd12195d1373bdaee874cb78eac8",
      x"23c2d158c6a5174ec493f2c05dfdec560cec9c794a0f247935e956fcdd7a7c6a",
      x"75e7874a559786bd9ad41ed623165a122de1ffbf8759259f4e644d22f1400065",
      x"8506338d10b6b0687154c1a5ba4af79033f8e132fa3682a3d9a08f99e45fbfc5",
      x"1056a0c35a32fa420a416a056277a4a37cc0ee4a93cde6a1815613cf79eec8a0",
      x"2b0c6c6cbccb5fc1c8888d5953a40a2803da87402bf782e558f4908f3986f369",
      x"90279cddf738f262257b1b83791fc3f389e5d14282e7a45f2c1a21ece2318afd",
      x"a490b634f86596595fc40184946216803682f40d4973a92ca579112ff5aac834",
      x"fd7fe233120ca3a3c52ef8d751f68f0e06adfe0443091d174c0eaf690453dc55",
      x"e5555927971987248129f74c02a17a6094a955c5295fbbc52c45d5f5adbbf216",
      x"1d50384fea4afdb80c658e5ace9bebae89641643e8c3ea6fc964ea827e7a7f0a",
      x"3720d0f7d38a96c896163f9752ee902e5f5ae4b1cdd648201532b78e4664c85a",
      x"67b560c2b2eb3aefab34e521ccd74ac8400eaa3eb4032eb3fed9feee21656623",
      x"fcba126992b6f351f9143a05deecc3ab7b1b5aa7285cab2d90251f81be63965c",
      x"56940a24ab723631b6a3648beeee63c8738b0b268b8564ec234388b2331967b1",
      x"381a30efdc6fe992733a7613324734d2266be41b8081531cdac0862ac8637b71",
      x"6d9676f424091057313dedd194b80e3b7ff067c9c57d50dbbf96ec65d436af98",
      x"75a281f5b85458e93d1031d6ec09985d0ce8fe793d73143a7e4210947ef776c5",
      x"afc96fc7bf1f773b0570b670dd64bde7d4294c9ebcf7571f2e0e47a68d4f2869",
      x"12fbfdc20f60824295bb61a3ed23da154116e1a312652e50d950f69aaf55e729",
      x"0fb4547a965148e7e467b870ba82f3ca8d526960abe6a097359587275d7dc0eb",
      x"ada63647036b150c006a9aa1ff5b94e2bdceb2b063c7c89752a8673e8dc43a29",
      x"dc03d9328c7ae534acdbb39832321c2dc54412adbbc8a9560d459bc9ea3ed3f1",
      x"32012c8988366d1f85b5e437d4a60bd7c428adfc3607a0d25852343f07f4fbf7",
      x"ef0b11501790472b313a42cc62d181f008dbd57826eeb4c823067893a7da203d",
      x"236940da9740095e7cd52c1cb3fbae8c497d980db9ea55f76da99477837bdedb",
      x"8636c2a965fdbe99b2c655ee9fea15dd344538713afa0114e587f5d1e502e236",
      x"ca2a55b394c79c39dbc4e896579b13ca0aff9a80602eba7d26938e7ab41729c8",
      x"9bafc100a1cf1e33b423f2565c90d839ddc47c21ec4c682ac4c37693888aae6d",
      x"0e8b9f518d2c62c3a4f5365e7a17d34e911261c7043a934ee411eec8b8d9a6da",
      x"85ba5ed2a7740c8e3b5ed1e1a4905592b606d73a2350e32e1b7e8f41de6f063b",
      x"92d68779b16c6b238a64c74a206ac7b92e90771e5927ffdccabc32c669ba751b",
      x"808fe7f620d5624405106e52f910b25c11aa34becd8bcf69ec40ff4e476da6c1",
      x"36e17b651d0278d46cac64fb8625de28b7a28f7c2bc8b5b243ee2765bbb244ef",
      x"f115548c82ac8adaf84673190e44aa6891a8c0f53dba21cdbdca9acdf34081aa",
      x"923099e53c9feebffa75b31a64f360a3516fd3e6fef481c91fca3d0f022be870",
      x"878f9706053bdfa34b22fe76a556e398b0cefcf4ba1fe69d84e165b831fde5c2",
      x"a0dd41ed8dab9dcac491656674f333ce5b0b32b19d6392d3fa45bef2bb6654b3",
      x"483d14afff56aede4b783616f2ef574c5210619a79aa368b61deb849d7b49ff0",
      x"166452f25d4730f275c05b0e0fda064d0fc1f3a79ace272917c2dba87aa6dd05",
      x"bb1a80af52265ea8057e01902589702fc0ea788478e1cfbb467636e6369fc1a9",
      x"353a43ac28bcd36995b00369bf9c6c9d909c275ff8c1a1b964881420edb728bf",
      x"7be8e6d695b122b88a0bd0901539a6cfcbc7731938cfad9a5e11e16c24fcce83",
      x"969cd0e8c832ed4c4fb2c4c1c96539a7a0d02af54e713754ef13a273bbdedcc0",
      x"9dbec61ab10420ec62f582bab065a87a6030b7753d65eaf8901a4e21f2b914d6",
      x"5e4615164ecde8e7732e8bd07ef6c3cc0f809aa3d8b73b98cafa391cd8723f5e",
      x"a6a6a164259ce35e8c495d818310a0e069ef39116516a4ecb15155456f644b70",
      x"9c5404e5c642f0a194217214f5ad57842239a9238d91bbc0d56f7df9eaf939c7",
      x"db5ebcdbca3c70d88fc36e4db39ab4315472a5f0b192aa6c614158e4d7aaab5d",
      x"bce8ddc0fb3efe0a6e6d32bd658025f676e0f03d0428566793aa5c4c5183666d",
      x"aa213e6c645b47c4b81969e7fb8da6ea5f865222292d974ca4e2eef8fdb3770d",
      x"4c31cc68d565200b10eb3b6ce69ff27e07a3b3d4f685149086176f49dfa7ec25",
      x"342aefcb8fbe2e82d734a47b6feec4316ca8bab5908f405997eb0fba1c2796e1",
      x"9479e57e065c3c4494ccdaef43f81733ee40b1021e86de5e027ddb49ea67d90f",
      x"c32e12a9468854e0357cf997e4fc24261935bd783ca8ff2f9255248edb3de45c",
      x"1b803a8f120e85dd715ad61e3355c64bf3bdf179c9a29284a62b89ef2c406918",
      x"c8dc5e97e6dce6e75743a4f1df9b755433228e12f6b8be26746f53bc4d238568",
      x"16971f7af82261f329f64ed731969e9932cf1ea57f6b092e52b1ffc35a0e652f",
      x"9ee90aa3de64cbf36b695ce4772f457c3269f3e3bc5f0e0016bb0b2fcea16aa2",
      x"c7d11324ec54ac8366ffc854db36a987e1d122fbfbe5b7a0a30df8660b01cf2d",
      x"1b2200808f1004824ea3f669538564797a39b71516c79c2f55c5849f9be6563e",
      x"1555301aa20c89845de0ad246aa16e0098bfb5ffaeee94a512ecdebc2e2c65e8",
      x"63214d7e181d2d81ff3229bcf5732c7178246f0435db48c67ef90db63310c3e9",
      x"3b9ebdca05e9853cdea074730e2c5761019a4ee010ae103ab49b3dc2a3152bb6",
      x"b7b365ed2aca2601a128858b459c93fa0ef0ed55018d0f743dcbf6e1a8e978ee",
      x"cec5a95c922d7613c2c0df1e98a16ab3b921a65498886300f6f116f88ef077e7",
      x"3f8468097db49c414aec3a2765f08166c96e7a71eb970662e8da63af558438f6",
      x"3aa5d84f9b067fe6399bb295703f75edeb20bdbd57406007979f6a6970742e52",
      x"0d5ee5db78f86a0d7d967093f415a550aadb61b24c600c9ecd2d4a14746f751f",
      x"a0938810be3ef1e506a1fec7845c31908e6b95281b1ce264d1210b0482b3e2a2",
      x"6be03530af1c6b89423e637598711f6cb8c1580d54b4c8aac12d8e87e52cec24",
      x"85d7b390daf24defb3bebf9a71fd0207988b040b30bed3b62cf8329191e72f1a",
      x"9d9da13107642160cbef6fa7a7e7e3fb5797b7ec307bf927d4cc09b5c1f83a60",
      x"9c073bbb8b4eaa91013967a853da08123061955cde89fd6407220008db9075d8",
      x"34040248e640a8cf180cc1997bf74433681666881158ec5c419e0c9854b073eb",
      x"523ff9073d4b54a14c3adf47ce1a1cadb67c4c87c99877dcc8b11fe77e65044e",
      x"cda698c2ade505c5051c85d895836e5bf957af65c200e4b97cb9a76e6dd70418",
      x"b2d22d0a19a5d5dd41145bb8a736e0397a77703f56bc977a9f7f095748138f3a",
      x"dccc702b2280beb39b61ae4a4b294828c615b663ffa1504e010c681edbe0bec6",
      x"976331fd67a0ce223c89c160c67ca785644466735f33b5d404b6b4ad8197a326",
      x"43d1d80cfaa12759efd167547a1e71996fe53c15d63e48bc6b31a6bb256f6749",
      x"70ffab37e0e2d246c7a2cf2065fcced4c13c630aca189cdc48a44a7c1367bc4f",
      x"db3f155d1580ff6935b7a43a0c1eed7fbb700b44883984ba3787b55f6d9f65be",
      x"7e14ef9b813b977709b880673384fbb139f47d4266556ad397d0af5cef9941c1",
      x"7283d40afa3ce13ea81769c74c4c5073a9b3c66817cb199572932590ef482c48",
      x"0a9d437837a165c125dc78e0b15b078a1708863cbf0aaaa56aad3b3ff64fcf72",
      x"8f163290ffb3085ffca0bdca0cff313dbf72a99964cdb205859fd86f882c4808",
      x"d13a0fba97e816d0fcfdd175944cb9fe5f3351cccda41b6d8794fe166032465f",
      x"81e62398b9fa05bdbad1bb65e63402fca081eb059ba32b68b7755c21cc0380f4",
      x"832b26778d91f22b422b3182fb24713f7c7f36405710a406e1944648b9250c45",
      x"e258e5ba06a7efe8bbcbfaa2a28e2b7d2343d3df17e9321cc8a7a6f039eefe97",
      x"26b158773a1b705bb6905f254bc39ac1b19805aae0a7bdb37a7a70a8557f249a",
      x"ac7460e45b481aa1ea0f6be4da6a2707734e846f9b630d4e4b4752753b8dd6db",
      x"ee5f50ce2485b7a39b819a10be423d08d68ba061b64b495c6c3b2878201fd4ef",
      x"0311811be498e526d32fe8e6c29c0b9fd3892ed4952bd2e5529f57680f0e1dfa",
      x"42d1f275ac663b30d993f5e278a6601b7a9885c905390f744e415a99f24615c2",
      x"a746b7b5e00d133e67f2ecb4da6dda7614ea63d413112f7cb863890cc2e26d1e",
      x"28f653fe850a1acce7df24b374ec70dcd83bc7f0e91297921902a31ac0d5fdf1",
      x"769b124177b101f52661b46c414819e0197355576a67becc4832d080f3d631e0",
      x"31ef98998ca254f7e7d551271caadb132232aadcc72de6a8e70d6c23778e70bf",
      x"1600ccea62dc1582d01980544210a302a6b105ce8d9bc36c26bf7522e13ef594",
      x"f0d9e6aa4fd7fe8a30efdb56127e195f8854e68df2c7328d5b868780c058d5d2",
      x"c19909f3c558531a4a6401a4ac08fab24f1405abe433d38e85095d57e8d7ca1c",
      x"269cc9cc8380758bb7fab3d247d5688577ad98a51793e2fa6c64ac8b8d6eff07",
      x"90c0a85513ff39e8691d548650efb7ca14568e4cf192650e06a294d2d6161e84",
      x"4b7127741bba0b465a829b2dcae0c21d4be8ef054fd2a6bb4bdf2d3ccb1a6c05",
      x"ec4346ba12c1842bc18a18e99eaa177cf34023331421711ed87237412d09a079",
      x"de953b5de5b1697bf92ae929198d5fc172fba8a097db1dbe76a1b7939fd94656",
      x"48c24e4cc62fc1df44bd9cc38d0effdd1e8e967240b572a9a78e449661180218",
      x"403f22c17b1a5b6b10ed380e8d4bc2f60d2da9e9bb8a0ca5c70dad3b99acd672",
      x"dbb2bb548252d77409f25a08113697c62d3d94236b34e01e0526eacef674a85e",
      x"f33aa6d8d2deb9ece3cc050777c56b847393ca4b4c725d5facd6def294c4b3ac",
      x"9d447a382c91c2119d2b08eb6e886bf487491609b96497856484211a578e84e0",
      x"4e10d2253ade17b2c56a5c91b0083d0e8b6ebee1bbceb683507fdd5bd2cdae86",
      x"9954d195c87baabacf84c0c32a04f48d1d5a7b4930e608fadabb1bf9d5e43ae2",
      x"cff3787079f35f3a4559a2cb7ac76e13c14f845a7e3a8ddc3c08bdd796fd395d",
      x"eee1626a3352dc48fee634c1006594e6733019ef5a7bd0ee7a256dc04c6107b6",
      x"0d26c1609793507126f417d7ce10da31a786bce98cf5dbd08991a1a89f9b1d4d",
      x"a0c8f290379d3c7213071b96249f6d863e48fe3dcfdccba5c7c560a327226b23",
      x"c679d54ef2e1c8779bc17246b98c706fea03173540c3aab2eb58416b4b705a83",
      x"f6988f910f049e19e30755407fa7f00587b06d44a193b7e0a74615de6e8b0e06",
      x"f9e4560daccf1ceb0095cfadef4fcfdaf0680c345c0765fcf4e9e9b0b9a5ebe2",
      x"1328f6ecb53933915dc2f71d3661652585f468aba8a92ca673c9de2817f2acad",
      x"160ec7372a172459c8aa6b07e2cb7c508d88d303d5036bd8fc059cae6555fd60",
      x"2027009947c0bbc8814bac46aef54ebeed2eb0954b0356b1e137846549305607",
      x"da662db328ddbed70c1ef4d09a5bb84b2ac288a5ec590a8947b198053c16d89d",
      x"6f058a035f2d98c630a40db33a2b4e07198536673dc0c7a0d6c006b267943915",
      x"b9791b427629f5208768d3e36a7bef1668ab0264d39386d8f6ece99872fa45d4",
      x"d75d14ba929c2b23e1c523f35f4d93c2e5b6fb6eae2f7f286a053df13235e144",
      x"77e2ba8acc39ba27fc707e191444c7f780a0f1ad2d543a15df53f2c22757149c",
      x"8ba15608e2fe20b191a9fe07979a51ffd19dbd8ba47b995ee24a9c73832e2e8a",
      x"9d11ffe65598239943c1536fa37fea29f14487b3b46cec73bb2fd07ca8ba7399",
      x"e1dbbbff33c1e2ea1d351827adc11d8f84760b03fd57c8b00dc7ab19f0d19d8d",
      x"1eaa7c17f338e7d413c70ba1194980d5e5beef4be27ed6cf7a1a4c9c3b70518f",
      x"65d71418f010093720667da972044f028a5ad131e5d117a7c0ed181389752611",
      x"b5d11cc7247f847e457f4271866aa29d48d1494ffd5d84484f2f675e231fca2e",
      x"794ce01f83459864d6354711da6a91ec5eb6488702eaac533ee2b28450b8edd0",
      x"5b6b94cf38b7e7acbe91036a7077b5c1bb14ee2e0f1aa67143645c8fc8005409",
      x"cac48e416cdd7e597341a78f097441295798afb68e4e3725743724c07205b3c7",
      x"148b89366d1195320e22f16720d361f0241a3bf1022c48033b4d0a4584af13a4",
      x"428dadad44023118c40b4268100c6f2abfa8ff80cc18e5d2219b2b398000c8ef",
      x"efd693d7e06b7fabfb440137f747841e6dd81362dc23b69281d9f662fc6a899d",
      x"5969d09ae9397c542f5f93572c0f1dba66f591beeec05d3a70600807de0de98d",
      x"3cb417f1707d25d36255676889f7c674294c7f5042841ee7dfef8e0525257804",
      x"a1da3bbe711f799b500d587e2dc6db2158e34dfc49e2246c489743e0fc17a011",
      x"d4c79c60192a90f0824a5bbb20efbb64a4bb2d381ea55c1a990c78bcfd0efcf4",
      x"c73d7b571c4aeec72409099365c50b8289db906a5d694a06c5735c83ece45a71",
      x"cce856dec4036ef1692523762ce6249043a41df9337174c40f624d5ddc616e9a",
      x"87dad393d0a7db74fba6b1f529fa434c7a7dfe26a6be1db33d9eb8b71dc36f80",
      x"d8e87d12b6f691e4c7dfe1cc6f6bbebed3d90a9701d5753962ca3a201a6b6851",
      x"f97dc135ba8605443d5ecfcf2cebcd416670c509fdba59ef7e8feba6c82a08a3",
      x"89dc4adc409291bb0c140fe3956d1318d04a5dc1eb5abc6fd00cd7f4a97d16cb",
      x"b014a2efdf8857871a8613215df68529fba588d0113444f5f36eb7ee33bb3f59",
      x"cdbc39aeb8bcae4282bb1a404baa9ab66fd978dee02f0f3dcc08f17d270030a3",
      x"ffdad451f9c0aa1700383e95a9127ae39b7c5c33b1b46f30c863453b4e23f2e5",
      x"d61e7af7b8141ff4cb2fc01e572e3b5ec72945b82e6b62c4e34336f90ffc3fe1",
      x"762d3bc15050ee9775bf94f57e9b7e3c0b4840ec16ea53ef024a967c94801e9f",
      x"550ce4cbee1f70ee75eeb83456a3591d80c0933e5e11e25054f1e08c9406140a",
      x"11256074b3854e3b8e4b363eb1098de6b3d5b3acf447b02f856c9814c21aa920",
      x"0346ae73ea83eba8302fac00e59c40b9e7a000742a0f4db30b694dc5a03f3c5f",
      x"5de6f76823a2986b875c916f0c8d625a77ca566be7d98b2ce8b47d293c00acee",
      x"20de125f6ef388c46fce2b67870b436fe2cf16c4ebaa2be858ca40d13d959f3d",
      x"061849881b73bd4c6dfef14297ed64f6bfa458d70305e5039120641e37076b84",
      x"d651ebed95b9c5258c196b4e64b7813930790eabb2921d11efc166fd514596fd",
      x"26e307f7b7426867c9c15b605fd5db13b4c65ce230e3a9aad798af76e3876e44",
      x"44f66eba5dc8e7fb3f478288c5e18ab3ca4bbb12a9a357a3b29564c634f4c629",
      x"c87ce84cbfaea957cb71ad981e5e3b75baf95d313ef7aa46012e0c893d003b93",
      x"5d8dd26666d3d6ace6a9f2184d3dd465e075b5cd11a482cd6ad1901d6f1124a2",
      x"28a27c605b1552e56b60db7a43c99532800247a90802ea0efa07aea2d32be4ed",
      x"4abbc2e1790b94aa732fb07906eca0959be757e9239a518de4498ca15c6d300d",
      x"8f85045c0ea7ef3d4c65cab44f420d884d47ad8b18c24abb6bfd22cc769686cd",
      x"9d2aad2ec7b88b8bf963c14fe7a731048f058fd57bfaa8b9f4d5810fd7421b9a",
      x"f2cc0d0528f3277471322155f4f504f4ed7a16018fd4248127985c59024a53b2",
      x"c5c76d28a7a0d657149bddd6e624d0f3b79e0c3b8d3e6b72a4e2eed58d893660",
      x"411d310c0785ebd37553cf381c65e22f412881974047f41d1b7df2eeed55dae6",
      x"1ffe7b997c17ec5dba89a3340f13458b60d79455ecfe07cc6cf09fd9888e5b20",
      x"0279eb19dca9cfe6fc4970773025d611a6f2ca71bdf25ae316ab63a5c0815a21",
      x"5888549db5c91658fce57e87e942f2f0776ff248d385c0d4b1d4b648425486c9",
      x"43c27d31ba4d2158034125b7f4c00b69c80d1f0c53c72b7ee793262259de829d",
      x"213605672652dc6e79e58e9a85aabe49f570a5f7f412f944aafe651b0195ae44",
      x"3399a7b63d466cd73db03ea3cf2d8bf6e9703301d51a86b0bcb5cbff1a12aa00"
    ),
    (
      x"6583f852c84d91de0de62afc6834eb6557446b4279abc5520614637e2b377198",
      x"1492ce9f89b6eaa3cfadea4a0040e5cb835915515464510a5c834b5d058038d5",
      x"49c09d1de5e23d2633640e8c97fd0982968c367c457667bbf7369c3cd822fd61",
      x"c0cddf0a9a1714c4595a5a77d84c6d0d4eee4b4792c84d2e3ed37cc46320b0df",
      x"db7b096d20ef68b2862cc19b16d4884062d021059289a3dbe4c01e9519837ffa",
      x"cd6bc6990c016d25fcc2093b6f55673a0dfaead995caf1143f6074d68b8be5ce",
      x"75b2e9916645189f20c5d3a6d80bcd24673dc6dbc1093f4eece18940701dcd00",
      x"82f2ac3d3aa80a11ecca4abc0abb721f19de63a96200dc0985faedbf236cec4a",
      x"e5a4f8210b637060c898bbc0caa652ef720b8143df5cc9f3576f48ba657d39d5",
      x"0b50a6d0798b9b0e584c8deb4c3855f9514cd959d571b21fc7758046a1d6280c",
      x"b4152345a900cb1dc2e711f390aca3b0af11e63145533b5945e9ab08acb30c4e",
      x"bb30c4510654f2256a3d03a981fd8e665d595ec9f03b7f2dae1fba58d2beb4c8",
      x"67eb10bed5e5d78c9fdd0ed0b0aad62a3fd1b99ce1bbffaaf32246d6b789c75d",
      x"7c26094440b3f90723e682cf9a0046b005940caca4f7bee44aebb172fb86d89f",
      x"c44291816ef97f0c9256dc7b97d1f1f043d518c498149fb3b4f300e10688eece",
      x"2e5fbc89911eedd27b751a202875dab8b970be62cc0c19d915e9471912bb66db",
      x"d62c17809f9fb3df56d3a22432c258898843f30dfc4f9507f23534faa84fa1f9",
      x"8f0aac7ad2abdaf23c95093f35dbc883cdda03e533bfadeca82092f0e722b05d",
      x"ad8a9106c4c19203749bb2f0fc5805e4646cbbb87f3201268fb4fee584be17d0",
      x"c5d9c51a4088953bef3ef4e37e656dd3abcd858d9c9f67efd5993aa859220205",
      x"1228cfa198657e9c6b237f6b6c044f6f230303a76d0f4589127706edba63e1e6",
      x"7af6571d2b4740331fc9709c0bc22355d4da217a85b355a386d5fda48a81a692",
      x"c4c483dabb0c3904106cc8150e59eab48d077398914c75f9d04c9072e4d4ceb1",
      x"720b3d098429ff99e8904892da85240e9104cbd4039f69cb7a8d00d648321979",
      x"ef97d65ed5b9634ff7e390939bcdc8c67339b30657e7e515d32a4c97bc69d1df",
      x"17fb1e3d3a122bc965d5614b70b58ee64c3a838769820caca84a2f3ed72d3a0b",
      x"eb2dce255260f230ffe6226d38e27d4676fbff34458c6735a3fa395526d9b4db",
      x"04a8858c78b21585d845d8e3c135d6751f2debce6d1f2aab124661d8432080f2",
      x"23e864c4f033e65425820b1bffa2045bb2bf740b9866530ff55b68c193e42226",
      x"6b031b41ec3f1f5981b4226842198ca24279791d1a80d677b1b759def19e7683",
      x"e829fb992ea9a856442b378e88813241d4dd93f8eb7267dee07d8f271aaac9ee",
      x"843208bb0e1aa1ca9fe20751e4132e9f0e90f143112969c093a97e1c58e755c1",
      x"d277fba6c5fc80467e4bf1147e3e24dbc6539d2cc8796982cc8fbac1bb6e3628",
      x"3b007df1a0139d881af8a20e82a2b6b52a49a23c1c8fd9a3fb8e489937063943",
      x"5075c51dc44faa7b2f460573ac0c0d4f7cac2ef81067c7b11f0bbb98f9c139bb",
      x"30260d6c659e6b9ea5e443767d0ecf1a25a35492ed9975490bb88660c29538be",
      x"1522f91481e5c37b7f17e01176a1736a392e33c9b8be64aac63e595b3a68accd",
      x"425a6d87428b184add4062e62445513af3f20f379e8b2f38ff27b5f4fad71145",
      x"588c700e85ee7d3f11ba07da4c6bdd61945d6d2fd9918b713ac83bbde834cae2",
      x"b85df4733fea88e45b4073d0e03de61ede7842a0b787acf60e9d2e05f188f8ab",
      x"e853069b3b5e15def45b8ea27d0d7a72948f8246f6ff0568f4fca8f25bdc55ff",
      x"ce0140ec6cd70a36e269b63dcb2250e4d15e4b0c235f3c866b13d94648ba6f89",
      x"22631f4030c96d28115e83c23bc9b356bbc446de5009e36e4ad62cf5ec5dcc3c",
      x"4808ea2f245287d15a1434e71713abd4d02ffc19d90a8de83b8819b2a3b5dff3",
      x"63bbe0e1e9efa729c556be2ee03bdd7df836fbc4ee82818787b84d8ae2874dbf",
      x"a7dd28d1268133644c65c56ad019e8294bee83ba4bbef903f48bd073294d3507",
      x"4f037005cdca5bc9c3f77d58128889be9dff1f68071dd26d7d2bfa4401a8d01b",
      x"cceaf83b193167fc80b3fe03ff20525bd9fe310c8ac5fe9ece784ba22d811548",
      x"2597413e488b9986dbf831ee46c1149b09244fac06a1fe2a67b758c0a4d1ad77",
      x"85534431b677f1405759355fe3d519d9dcf95ad5c665c3710d1226e916205409",
      x"51533c9522c94b4b90503d91f9fce0002206c0cec54781d58127fecb0dd9f1fc",
      x"7fc1746096ec0f8ab240f20f3812e2db5eb9e14164062ff00cd5e1a4ddb7caaf",
      x"6dcef8a5a312864b255f81151db27039077f0d217f07ef16f48d4dd3b3fb7226",
      x"500231e93e045ed6e708609a8f01a9148e3b93835bed60a4e363544463b8fe01",
      x"42b6bd7933d33c19061c5bfda3ccdb4d49613d18abaa9ab79a3b0195788796cb",
      x"838de61c5a4a83943f3ec93c2bf04e988928486cb795f9610b66202f9ae1f804",
      x"6270849cdabcda6f4fbf1b3891e422f37677dd74d2dda05f647b59ee6324d9ca",
      x"69ecf393c1ecb93910308bae839e4fa118b2bffed30a554cb13392727c192858",
      x"cc73970c50292b75e93114c0c27cbd4e685b9e4decec3f43e7a09a4e5526e0a1",
      x"51de1418cad5433ee950fa4e2e13eae706c1ecdee54342e4b147cbbc2ca99749",
      x"312412dfec22cb455be2ae7796c365d8e8ea4618e204e49efccd0538e1ca8b3a",
      x"8d2c9795fc50cf93544a46f71061c6c24bea01b6c1929c0ffc83de4b7fb6ba3b",
      x"13e135de5673db57e610827c8eeb2f926001b11f0d01d82f1ac8bdfac0f96d4d",
      x"4a8ff0ca51dddf83c5d411fef5d1bda90f7e88d819ac3016d92e741fb9381218",
      x"039b9e907630a47ae6926bd429582769ea2e0ad2837e040d0f795dd41e56a58c",
      x"3e1074f3566d36374f6afd8fb233817434ca2b19cd6f2c4f7387885ca3edd5fd",
      x"7262da7618e58c81bd8f9d76cabb508d74c07cf018e6ebb7b5bdfe85f46d0351",
      x"2e4346c4b80a3da49188b54cb1a17106f58b866e96e1045106e5754aa000f38e",
      x"f4cdd6c627b82014bfd1a3a144c7a677f387a0a0c957354095bf9105116661b1",
      x"83e75fb7c49444491cf4e44670b84483e1809397bcd9b2771ed2987647900c7a",
      x"a1f99602b9bcf2de9e3f4ab7b6c5bbcc492c6f1ae1f7bf1b52d5ec3056f515b8",
      x"817347922e24de5a03764444635137363204edbca3ae32e18e3067cfdd51d5a8",
      x"cb57165fb28e7f468daeb4bb2e014ac5ab7f72419ec0ff1c43ca3cad48f5a913",
      x"5fe40ccbb3d80b75e5eee0e670e6ddf6ecb92dec13d2a6e7fb94e6ad9430c325",
      x"7de4dd5513a1c306fd26e6077551526b3e1fba9c07d2c741c2acc0e667409be8",
      x"542e796962142b9b02239776bcb9f69532708a062dd446ca6ccf0086c0e7bf30",
      x"7feda1b0608d9688c7a2da583864f1882e54fe9afc04f5de78b9e60dd96002c4",
      x"882821b63feb22dbe7761e9655f5feb2851fd04847ec50955ce73de631a70dde",
      x"f7164fad7056aff99c212d79c334f0b52f55f6a973fbd0d8b2441b8f4c886319",
      x"70ddcee7fdaaf6ed5e07606b92232e428d02de9e0faa9fbf3173ae336cbb7413",
      x"42e5759b585273005119b1006489bdc7376279615413d2d40a37efb17bdabf99",
      x"e1fc312af1e33fa9c9c01270843ad3d4e02b87d17873e07607d12ea609fa3821",
      x"69294cf6da4e888e53a30451bb6ea2dae54ea32da6166f47f4e96e4b50c6936b",
      x"a91783aefb95ddf6aff20906772046d3108c590346c258b22cbf45dd5c4e853c",
      x"4db6a92a8c3d5ff0c8c5819f4fefa859f134f263b85e02db3e8df3f445f7aa73",
      x"d9891304853b9d2e6a2d63d58e567c3aab42e571c9713f48c6eb8f2dc1be0e5b",
      x"84d865e93d0e0ba6ab0163bf2d4a18b68ad29cba77b09a6c2f10d6e4b0afb994",
      x"8aa28a173ab9116647feb235a5251a80211119efb78cee04136385bbcdf4f438",
      x"1f11b5f6b9f2a3933b6dae32f51016e861cbd817f19e94eedab580c6a573b285",
      x"7ca562c625dbe63c0607bddf1c3cb1d5fdbdb7683184b1e72d1bed045898f252",
      x"cad1c3acebce56db0139c786498198c6655308951361f4ef1963f30c841e117b",
      x"b69a3892757143fb5a2905eda5c41ae44a4f38bef80fd64b5d2f94bb526d377e",
      x"4b094063d70b4f162a538211b1c664bd5eadd7c65e607561c866599b9ee5676e",
      x"08f7daf65ba8d28acc5a8f18f97bb9b66d5da39cd209e8a74ec504a59f51072a",
      x"508b8464eb46fcb79f1074a1e9610a6eb8b5c97aa1c2656397064be4a89cf902",
      x"5e8d8cad10ed45659c49db7f6770aa5655aeb8235d26936d4f381f903e0d9250",
      x"614f8f8f8474a35033c57cbce93f7e70d17b32a91ccf23c2f587cd7bf13a5d17",
      x"218141323943c6244deeddc021cd39c31173bf8badc5f88894160fad04c35f7a",
      x"96966b95ca7550851a768b1835606d5a6ed05e120187e3d1b11abd5681544224",
      x"3b4b8e9159306ab49dbc00affa16efc6a0b03c452a44e4623348e4b4c54cdb52",
      x"66997efcd148350455f83c987cbd508922914e74959291b032a6023364d17a33",
      x"3b3c1d02cb4e5f4ea855a9c274d6cd066e4b7e2dc97bb6b4e859a7f2c1913ec6",
      x"e3e2f757f1d54451271daec27326f54be50ae744a9ec6cd565e3dd3cf65749d4",
      x"df096cc1b1af5462aa4dbd38041f3600c9218a10e30252ae31556e3eb819adb4",
      x"f161d6d7ca52c31f0643100d233fe1bd87f6c5bb7fbf8e5a5f86837c21b46e61",
      x"72178e79a92cca1fddd415cc29ebc53c9c6d16518495a3dfec50b7b99a99684f",
      x"7b1e36aa215b407a06b8e1b92ad93ea48521aa8299b7d8cf19952d9b0daa7fdc",
      x"6629474dbb69ad6b6c11972c9562eac03a30632281e5974f673297eb1c1abd22",
      x"52276ea3de456ce438d2f2328e859235edb0670ce01e074a73ba64b4656d22e2",
      x"715eeb18dde95a2491a7eea2f9d7ee4c839e1a0a202a123b0a6fcb32812e33aa",
      x"a5f5e618e0a122d957a623a73ff4eed02b640b6f9138d7b50ebe48dd0aad2dd8",
      x"34d919119c46aac38334824b408aee2e50a19da24148a1ec4b5ce50640d9a0d6",
      x"c58b8589ddb93fa133722ab6e402bb5bd0782dde7ed9ce384ea946cba7252543",
      x"95c0f013ba0d0ea90bd8cce260ea60bec25e7e4f4fdb1ee7511e356252c232b3",
      x"ef2d30cb73cdf3dd95cb6778241006e34188bf372e8ea9c518f47bc29afcb768",
      x"6f5fd261b0071316d8a462e90dbc9ef6c198137a869f7d79d38602c7fccfacec",
      x"1983dda6af9f7c8bd2d0ec20beb6f578f9614ca3691c6858ab16cd8b6301e0e2",
      x"f4efea31c04345ef3550fd6ea5aa81e89c13f814bbe078c642fb73bd0f458f58",
      x"c170783803b8c3b31844bf876a42f78e3ea7c69693ef2b8ca232cce978602be1",
      x"6737d4836a7a7a69d817f340fe3cbc377073b00d34ec05ce73c80a04e2e63943",
      x"c38fd15a414021ac159fa4d3964e6becd7feddbf56d5cfc613bcb32cac774678",
      x"99db06235f403220a5e92d105ed6dbea803bdc5fcef80717e19f57f45bd1d82a",
      x"9757c4acdd32b5b462c62a4f1844248afbcebd82754303eb9f008a07cbb24c4c",
      x"82c17ae19707a9ef78ff6f98f04eb6e6ba0ab45ec98231f181e9aaf478b18b98",
      x"387c0d8fa0e2cef122e09e30119065982e3ff5f8f37fce233e283626ad042db9",
      x"8e9bc707528742aa58deecc257193356b6644a5ab25a2475ac59dd143e335586",
      x"d47bc505e3223e07c6bbe6372a36db84f11fcd6748d05cc77a6e18bb8af19e87",
      x"ffd472ad97bc336609ccde97477d47c39cb51f8f0559d40829bf904674555ea4",
      x"a52032681468eb154f9a7bcd12877e923a0c03fbf195d60017a6139633a22101",
      x"3f766f6261e17f96b89ae2dbbb203dcde7e7279f7e62faf5000bfd4de774e05f",
      x"b4e74580cfecd04af5172cc29206ee30bab6a3cda583094a1c33644f2260edad",
      x"c82224bcb10ed83cc4b82ca5b2f6a57170163e8f81ab9fda31528884bd6b7cbe",
      x"9ad8b159a2b43a435aec80d8e1d73cecfb6ae6acd658005d722f918a54937352",
      x"77842a8d0231a22c1b3c24d1129bbadbffcec891baa134008c8f59f08829b64b",
      x"fc22baa781b51d2165ad5d6da79362c5d2cdaecdbb404569554edcdc7272baae",
      x"d0ae05e8df5f9cdcbe95e59e30cd8573f622ead991f2d1a6654518ae0ecc3c0d",
      x"03bb9b54fda258d46dc1c16ba8537923284f78d1fe42c9c08eedf1523a183595",
      x"e4bfb3f5d457619c185b1ec6b77d855c543c96c03bee1bf6c1cc0b08e18d8654",
      x"11d62fce862bf7d9fef97b5d468b9f0f845ad6196c7ed952fbf90930eb71e2f3",
      x"d01c9d365937b728da793ba1c2621e6eea6bba039556538fc1b0821d37992cff",
      x"5f8b417755ae74491d6cadd9753a0425312c91ec9f970d090dff167d996585fc",
      x"37e370efe5671deac03d094065ae768165a4296518d0d6541a8e0b1f7924b53e",
      x"50761a9385f890a769a6e4ed50b00b0d987003a785ee378d9feb5609c162a8c6",
      x"8653a71cd58f220670c24d32056085d589dd153a1d55576761a415cc1c729736",
      x"2ae50b158740e1a68398c24e2961b3757426618d790f55803eaf5fa036b7e2a1",
      x"5b5b4f2d3b444cf28b217837afd2390c9355cdcc6fb2b29e84e0fe6b324caf2d",
      x"67e6b4abaee7974ef6581d3b8e10c74f2d0018820deee486c8ea1dbb76a33344",
      x"1d446f696e553e6cc1907e9bb3532dbcd6643bf1eb55a17b40f34b8f474a565a",
      x"89c3997dd53a17feac08540aa6ea21b54b82c7accf75507594f36a4fd448bf12",
      x"c04188c083345741125fabbc1cd4ebacaa84aedd4819ed53ee0f94e7efcb2f01",
      x"5ae7f0f6616991a4555259571a2bb71ba29667e143aad5070901fec7a51ff4a3",
      x"7f6be56e0e4d3bb4f7cf2a0bf0b7b5bb51414536a44fa2b764a8ad095875b51a",
      x"94234f1482e6079299d7fe4fd3e9447b12eb48ade48997a875c8b131f7fe888b",
      x"1143bfa697e281113c2b12d274eb02c5cfc4d6accee0b9d70b9e64849cbb25e3",
      x"12c0d6b351665468adc8f924e11fa7f591d30535b15b20009a47f3a3af0dc213",
      x"32772f98103b5fd8f50baac92f597cbb7ecb8007207d7b33aa38ae31676b56d5",
      x"374308206f4a7f7a0aa67e1f73a8c64298348b6e94ac7501b8284fb4fbb02cf2",
      x"3a33a88c6bd54ad331291ac4a2b5bd894233d82f0dd395633ae90935d2b51b61",
      x"1dc50c274b4b7dd85aca29233f829b224a7352863f18da137ef52610ae7f6f74",
      x"64551e7415020286d3ca31cf1b23c64173666b3c17087da42bcf5748b23c59a2",
      x"b745c5b512efc81ea5af3aa88ff6aa4b4fc394d8b3120a9e3a05cf81d8a6220e",
      x"c87d03eac0e1cab4e031f8da48a9e3e28d3c59374a5d15ee2b69542f44e05e69",
      x"5dc099818a00294395d5d9c52d31b3da6be28edf36dbcaf1aa310ad235523f46",
      x"2e19a4a3abf73ccd5f59f41c5c543255cd644f93139cc31899c195a5c3d88e2c",
      x"43422a9d94d549bb2b1183f0701ed39d59de89a201b5a2b34100753fae18fd9e",
      x"03635b4319108d16102046aa92e2a3edacf1388888401243d976db6554863cbd",
      x"eaf8a23bf8c10fed353eb4313cf6ee0c59bc4bc9b7f7d81ce871a230c5610a56",
      x"bc4873ea251c6c93b2aad50d30eae2eacc18634ff1b33a77f9e038e4a2579a3a",
      x"417fe841c5e14bb3c8b40bd94e7966e2477009bf2ca9b45300612d57d830339c",
      x"7bef0c63ff4065dfd624259d1183944c1cd1f3fd85e38d8a9d75e6ed87901cd8",
      x"db6d4757765064889a8405133cdd3fc73f9a1fb0d401e0487cc5889ab014aab5",
      x"6abaeed1ac0e7cbed9ec2ff5bd53a06ed28fd9cdd9d7d8a8d87238cbb1709ec7",
      x"f27f9a02abb32e8bb8df57dad6ce44aff8707e23eb86dce36c903d67c5e4a0e8",
      x"b525001636eefa7f596641087215f73db99a13072f02d9c72a6a358e7584c0e0",
      x"004c3e5c4b0aaca1d06d3d94a9b86cdd7edb521dcf86227851e84f5b4c7325b9",
      x"274bdcf6314b5213863f403875db82380dc820af9ad9d767fc16a4dc0c2112c1",
      x"95f060878cd569cbf68adb6eefd747db25afcdd37eccf809aa0badbda28b42bf",
      x"a10e199f31541dd4035b6290b6c74f5bb294687eff4e82ed0e1b3b428936a1b8",
      x"08b910b27040feee0b4c5705199c0933d3948c5dffed877327c2522b75118a41",
      x"51374568c906f02e45637d3e322dc975ca9cc04b18f17f25332d270a2319498d",
      x"8bce904bd11e7d298f38da5f691ba37224233f822aa98e4e18fe8a289b1ee851",
      x"56cce305f56b2db792a62b5517671abef2e9e46053d910b61b2e9453d5809bc3",
      x"cefcecd8288f7230c59fdc0ecf51a9b65ff38e3b71f9d4e0cd27e17c0d5c0229",
      x"2224790dde8d27c26da33ae05f2e80d739e9761cd574507e83f5374aac84143b",
      x"a6d7c218956768087780b4a0843766fb09caa0509fc1e9e936a9040b8b177fcb",
      x"e4627b8dfccabd510c281570fbf7cd94d6bc6e755800601b6b733acde38f8671",
      x"6f6563d0a45e5dfa2637c48a4bf72ef0b7a71dd1ade9583b6cbb8c586c6a99f5",
      x"450053d1970000dc2754b7a6416b7df0d42578c9582c770a35801529dd0e8215",
      x"96f441a909b89abdcfea8e39fcbda82773cfaf57db47d3b7a6eea69056fa4f4b",
      x"639679cd33a39e6f6902019ce9112ea4501b53ed4f70dbfe02a14fe94f3dff6c",
      x"cec36c651249f653fecc47c41c65850d95b54ba6a5a038728dfa4b7d0476d695",
      x"69baa0e2e3fc8340e613f0ee115ebad03b00ffe14ad20fe879a14da5e5828bd8",
      x"7c347af474d3b050644d7596e9bc84d2b7cc6f5f090dff44ce6842efa1326b10",
      x"ef5ca7e2135f084283bb98798567814654d4881d1fdbef3b30346757e0d2bf10",
      x"2af041b47b668340cdbb2515ddcc2bd575a84230f945b4704cde93aaaccb3b17",
      x"2d8b939a7a8258bb933a186e98e7c1de842f061da9ffc8252f03ce7a6ffc734b",
      x"76a580690fa24456f37b40a51188f037dbde6f29ee2de1f3b52625bc8fdbcee1",
      x"802317262107e37d4137e9cf9206ea91cf09a7ff7d11882522b6895a511a621c",
      x"44e2347bea8312ae1965cc9aa7b80e1473709cd465aca8f41f590a8b1e66ae79",
      x"3631d94badee522945aaef9b2c30329efc84c9270b2ad80c10cb0378ad2a16f0",
      x"ca150184c2c4adb11f0ee78c37adda1d427c67836b4b2f1826fb5a388d8dfdd6",
      x"d8c41023bf55263faca6e4c5484de01a16e81e92d70bde260755560dbfc8aea0",
      x"365e8c3982135a4c1e8a1302bdb1ed78948d31e5c40b3c118b9cb46cc542f266",
      x"06b9568e0fbe1b036f51b037f869898c8017bd46ce7a20415caf9149b584f066",
      x"a3ce8048a12bdc1e38b801947e6d4d14a7d364d33857266e1bb7134d2d4f2ce7",
      x"0f2dc7eaf3dd7c81b5568762fa23274a7ccb4aa3320f2b67eda3ae7ef9703dac",
      x"aa1bce951bc4bd1c69a7f3dd119d85ffb15dc2e699b49925911a47eda20841f9",
      x"d2a12c01b4666e93139f99fc1d60747b2fb6bd2b1c9dbe29af516583cf140efc",
      x"4b2e2274ce37ef4a9f0ecc71dc247af305dba672a958e641b720636b4235ff51",
      x"b76f0e5a8cc07bed1c8f67a532b0b9d0ad1a2380c3fa821321cc54f823b60121",
      x"d9f930e14b42d2ec5bbc5438230c3d6c577a709c672c0bd43542d333b145d1ee",
      x"93b4a09bbf3f186e51a4ed52b4365d7ba33d9edfa126e16a1a9566256b998102",
      x"2a07f433070e93576ddd088a70f6a71bb8deee0896c072d868473d566cb82eb0",
      x"7e6b75f73d48584677cc45bafbd35d629f3db79f5fd97ef11eb6e8fa7a0de992",
      x"e289d723980bb817bcddf9c5edc48f568329eb07650b6ebd575843a7e0b7f086",
      x"e88ebbb2461c6a97b14af22a99de9747538d717b9f56b7633fcea0b417e1ae48",
      x"79a7c1653993b3833ac14ecddf464485fd5dc6f7482b635a23fa811e42e4ee40",
      x"caa63aefd9c9e0d812eae6614dc731e74ba5d529087a4ad7e995a00c236f2684",
      x"9b949324c27a3261054c2d357d242e235abef5431e599ea2e6b29a9b80129cda",
      x"06162d5a34b5b9e5b758d8484b546476fd93f01f42439615b8724e99c1318ef1",
      x"21e81ab1eba73e617ed098d8b67f37d300e345b6db9489970d3da403a493900b",
      x"1a82642db7686a64b76613ea09cfcbd38c11e33e0aead4d7471b1e0887787d19",
      x"c840dabf915e51a1b8f28c6bbc0c32f95705ad0cb8af9f13e4f6c8f10547af72",
      x"18953e4f29491471f558a2c0326eca9f6056524a45d6a533b2394c646ad15430",
      x"78aae5f888cc206e5d1dd0b03fc59a22dfc1ddf5860d54a808624e2e1a35fff8",
      x"7b07c7e82fb96bba7e7ae5c96ea70cfcd2f51a31650cc647016029f10a6e637c",
      x"b7867a6d8ae60f16b42220d1ec13f6c427476d5a0caa07d8d8fb0de2d1ba7659",
      x"c3257cbbf43e962e8810843becb905fbf3b726d54993bdcaec7ddc7dea6d2cad",
      x"6388caa8676fbcd95fbfa11b33145669845ee4025240a83329dfa2072e36ea51",
      x"ee6d1771548e7a5b5ed9ff8043e68906a7fa222958a0b7be71f3e32100e59986",
      x"5f49cabe877b439225c762d4692ca89f4f01bb209e2ea2591b1ab2def8d33090",
      x"ae43f138d85aa16f0e08041944b3e1ac54aead31b39bdfb66f8fec16b8368525",
      x"481f2862d0370ee5d6ab6774f24e054c534a3e6205713aadbdb3175a18c0c041",
      x"98f862973e88aa064c51e91c0882c65c2d3981b9e6f47d8575d0931d69c63fb8",
      x"5600f5b6cbcd4d28603dca3cb7a042e70f4d6b54dc7959697569db685228fc5f",
      x"60ed538b2b0bb794b5911fb0a5373abdfa5d9857e18ea04254bf641a8c54c3a2",
      x"202ef33d93e7a1bb63872b0cdb79a7464c5bf640c5014a87636aef92edd8b6af",
      x"442863a2b022f6663632055c355337a69e9ca3bbe6c0d99b7378a49a7478c39e",
      x"23e953f21aaad130ea51e0ade67b7d838738be2f7004d5963c9ed4c9b3ff9ca1",
      x"007cce6ed8ee14f05e04555f4419b7f26fccdc2cf5dfcf91ca0b3a408c6e2ac5",
      x"d9864b48a64e3a665829b32ce57d7d323ddd927d5e0bb928f0977c88615d4f85",
      x"8e2545367c595f27a640fcf0451437985d493baba06015b49befaa155a7e1a5b",
      x"65ed179d1c87f7260b8dd95244c9202310de728bb302a15020f6b344b1d1f5dc",
      x"bc9a389f8631deced7465cfe2c1ac3363868692ae4dd510abdac45908c400848",
      x"0a7f708e61318c4021dd6cdf2ba42463e02ddc482a2f8c106c6bfbff86b48526",
      x"cff76ecaf2dc4ed5dd08e71d72e2bae3924db27cfd4d6d3074765e9880150b2e",
      x"c4b43c1d22bacb0205563f6accc3f0ab2ac28b2741497060b45f5471484f3d70",
      x"a4f6a507068c7567093f7ec300ed7e4c89359febc36b21687c4a157d53a2d28c",
      x"252f4e98b62262db8187b94a76a5cb6b79f23bc2c8a521de3a14fc2c9bbbf5b5",
      x"e63a067a4cb640a387357426f4986a8e42e90a47b8576bc7c19c36a517d25b05",
      x"b93ff6982a03c22aef56247b30f7f39efb8cf34e356109bfdfe5a7534702cbb4",
      x"10f497f4ef68f4af3cd326ad76ffb906cc85e7fb0cd79da5a27b49e05d4bf4d7",
      x"1b3ff8a00c62b4873a336acb6818740438098c6284ebd04483556b8f6b80be5c",
      x"eea82615941c8fbe6cd6070c508049e94f2fa3d8e2b8c0623d8161a33ed1124c",
      x"8a06c4ed7afa2b6ae63446b8fa340e402b24407359a3499889b2814f90abca95",
      x"29222bacb94d97fa565b07a30ae44ad89855cd941ec914aaf36a1451d5021516"
    ),
    (
      x"06e909aeac07597964a2748866e4326443458776acdcfa04055a0bb4855c2e56",
      x"6a97588c48666b56a7ffd0f07895b3e655806d29dfb22d1c57db1379b4ec061a",
      x"86c53ead99903ef47e4d645a87dbfb0c56e0ec87a67104cb764ea7fef9e9a12d",
      x"29a1c86277e11b8f4e9d96cc1140721188e4034173a168354ce63c906e7e9b66",
      x"f546dfe73e708fe3533882ba33417adfcd1933f9bd07078440a0af6ce420a3de",
      x"11727dfade493b0b358e68897bbd53df2a07fd9c6ba65ecfcc4b852eacff1e0e",
      x"b4aa5d124b3651679c78bdff04af856eaa74b9d0d91d2c38c8b4e2b0c9bde69c",
      x"7abff3a5c7ae3b09ccbb89895d252544101c14464331dd1d5b6b9a3628c50da8",
      x"4d43a1d5cafa40bdd044da2d37fe1e5e318f8ea112fdff33d78179faef64ef8a",
      x"38901e59845aba2eb8c25ec78ea625b82625810ade1d834b39a20e8eea2ca701",
      x"3b5d72795d5bac708439d83639628334077da4af79e2035f6d879ac744e53fba",
      x"06af56dd3892cd05c132beeaf7c06cbe0cc24d0c2a269004f6725d029d9b3e92",
      x"c1b5e59946286afa815d56959bba8bb6a9e4e0269f2ce560938b5c016b11a281",
      x"2203ae6dddf15b6aaa42e1ce2ba05241187176ddf2ef5f3880d54bd4d92cc363",
      x"7f443c9580d767050e21540bd0c016991b270663608698b2e813161d0d33efd5",
      x"c9e376aff5599e020d040e81ce5974f45bbf59be28bce0aa28fa22e1b7c64328",
      x"815d2c742ad6972beb8d648f1ebfcaff74e176cc4cc3e7cc5c081de2afa004ab",
      x"7ad05fb2b9cc410d4f22f6aa2b538bd5bc4074cb1cbe928f43663908d1ef8e72",
      x"27932fd65ad9852e4afdaa8a15f41bd56aa153af446d2ce3a92a28b4e24dd0e6",
      x"a251f3c45b4bc2127cd5e1a908702fd06eb943209a31fc45813943740b1e09f2",
      x"6fdd7e2cd4e4a78963596a47aa29a1c314a1b21cec304d097d39cd5f28c94e11",
      x"4042b0e132d5f841b094b7c399902e087b9890469f233d70ea4a59dc618495c9",
      x"e1483b13787fb9a99794cd70b06e941729b711fca79be8113b3c0ce5747ca47c",
      x"f13ca970c1a8a200df7506baca05d33add40710496251b1c92b01fa692eb16e9",
      x"af63001d4350044e91520e56e36e8901eb3de15bfa4523bdf69456ecbe57e420",
      x"58fef8e68f00b4442521ee77b9bd55ffd8d0e3b3f3e9f5c773c174132d8925ad",
      x"be8e0a6297086188152b7adddcf8c8deb683c8131d4015d8c9c9c76b812d3955",
      x"09823c3a5d712ea90d905a4aa4f96709e2c94c173a1cc7a2faa13e6fdb81fe31",
      x"1853df99c07df8369c96046e25e8dd9f40b96f714ad0be7bd674ab27f2bbc477",
      x"499f96395ac27825d16d8f307a586c17f2fc764788ddefa34518bdbde7ac49c2",
      x"a4af03467cf6c3cbb4fc329d9022ea8a60f05bb7c49acb01ebe00f8e122bd1c5",
      x"5b7632091109d720f42df4a65fc518a85d38d472024ecf39222e67d355c3f651",
      x"ec869b371c4a150098298f49885c42bf7387c958ddd9d254a65c3fa1521edde0",
      x"2ac9f9d9b8ba8437f5a6ca4f57ec98d78cd1e5fb13da40a7bba6d92cda803d9b",
      x"235afbf35afb1cfee927fbc91c83a8d9a47ecdd10151110b94a448e90a558b53",
      x"bc8929a9983b38865f6e3c1716adfa8f44a9f45d2ab97c70cf069722527ab628",
      x"f4fdf693584dd59d9ad0588c05852e6803b89494073b566f78e97515df131872",
      x"a166fc791a3742820de1edcb103e7f625a0dfa82bab6e3b1f2f04d58f8d44e09",
      x"a2bf95ab507700e0c16a5a2eb5dc8dcf08e72fefc0bd6f9fd3014b1842b158c5",
      x"4206c2dd785c18522fa6df01bae093849f185f9842bf0aca8d971e8e3c471823",
      x"42ff370d1d3ebe85b336782eacb10a505cd06518ae528ec964ea612f459d955a",
      x"183bf726988f24db879e41ad64e2330697388c5a8f5f2cb894a1e6880acd0ff2",
      x"9b53372cdbfb65a227bd21f62d397361889918cfc9c587da8a567b6c5adbe6f3",
      x"f61f9ec4436db19263a9ba520338533cebbc5c07754e0a8b0b66046902a530fa",
      x"7134ded9353e00654f103123acef9a949daeb0d77de8e2f68e01c129330debcf",
      x"fa0a5efd03681818b1694c40ab961858389970e0c830fd33c56ca85164ebde24",
      x"a3fd5543539d3190d1c7acb549e5a544775850b4626ae11fb6c429d0e9658dc0",
      x"3c6ab58809b91c01579464411709593947063284a4d42be9624f66ffbe489b6a",
      x"bdf0e3c2aafe7109273f2232c6b6196cb3bc18cc6de4a663c06413b792c12f61",
      x"0b073139a8cefe7ea3bf8d2272b30bca34c67d82916ab619ec07b0399f939d02",
      x"f4309d745bcd8203eb9025aff4d2b26e1d7ecc258bbd315c40eb620249b84155",
      x"4079fad1662cbf12bd12af505a5cbbdee6cf1f4da50ba4b54dde164f0756e358",
      x"686c2d9b6e801544a460b3b6b6bcb6232dae1a993aae02af05e6a0f1e374a7d2",
      x"449d0f596b644118b1ce8f1bff70bafc7afab206c1bf7c2566df6eedaa4a47d3",
      x"c0657d22b4940208f6e2fbc452625e17e433b4618bc5353537e2fc033bf0b721",
      x"1b95bba074b11048d8d848303d2de6158eb2938e74f9665691ca974cefc9f007",
      x"6bcc2be33b61ff82f0e7d8ab8bf44cacbbd8a2224dfde152d829fbc879c6e4ac",
      x"9b5ea8a7b3aa2031e460517b7df4883585aa81d9d2df82bcab0a7a00aa134850",
      x"e6655dddf3dab803017ee744de88889116c9734d0451c079272d17a5d6794e0b",
      x"42837266e84c27c5c0d4427d410ae35e006a24dfcd1ec8f893266bf0a8a04169",
      x"8e9e85e10878e9c5efd6b617ffc98198241f9efcf202b303f5238e84805519da",
      x"6d9a586fe8e2f65335022572ec77ad01b349cffa9fe415fcffe7841eae76c738",
      x"ad872ff383dca939668256863e9bd93bc345f7bee4e3dba522d07c21f36a6d89",
      x"20fbe14f1df9fda01e94b6918ad7b4241d04bfd7f1ea9f30bb5d4fbd3b930373",
      x"12e2a53be041c6dc103913994c66355c25b0f5ffdd02dda6d3aadad1a22b4e8b",
      x"719eb01f3bb7d90c7a54684525c6caa68ba19a52f83665d27484ce7e6da59497",
      x"37db1ec250eab6d9d10c6746f7f91a6ac6340639926d6d77fa647f0d5ecb8385",
      x"050a6d99daa5813d2b2c64ae68357f900fd641f3659d8da057cee08eb2803db9",
      x"0ed11f808839d03ab9798a544e232891203fcc24233fb521e61d0f854f9ca5a6",
      x"fd7ff7b2a0df81918cf969ef2d1a487d9e5faae6f4e39849524d4339eef31cd4",
      x"38c5292c6398de117a6532fb33c978d2461c32543875bf2c6253965b01944ab7",
      x"c649d9c8f6de0384c2b3b445229cc6ed29a1747d678c25a1d9460dec56170231",
      x"44e10c25a75adb3646440eb31d3f2d3e307a4d26c20d483d58c7f437b06c6d84",
      x"dbc39ee9e18083749fcdfcbffae9f93fe28e87f0a2c6670a7cafcefc26139522",
      x"aeda9e7e026ae02dcbf286b10e8467eeff051fc75b6931db9ceeafa847df30bc",
      x"b9cd16ded6ec4f87316df04005139ab4827de9a9b53f85f457e5dbbfe3e85c5b",
      x"c8720ebb23c8df977a2a076fec52196dffdddcecb6a1981ed34e296aca44d723",
      x"ddaf901443a0762223f94d90989a80e45fd98bd5bfce4eef489b3809bf14e0dd",
      x"8a3da3cb0c1a6d39625f96d5b9404e94808d841cd9ece55e9ea515133f5e5478",
      x"cb332acbe47cb126ad3a57f592345ac953a7483e25771c9d82a3e534a1979d33",
      x"3c42d3be3aa66d47ff4cfa857e47dcfba378cc6e8c18206186f6e0aeadfe9255",
      x"1aa6a32bb01a84f48bb72f78821d7112077e3e07de2171dab3ada625b8bab807",
      x"af606d72a512f8918a1c7dbff8153acac3fbe1992ad1b7f67064b788b4ddcf84",
      x"f47b591d6051aa89b75bb5e131707ea11187f1568959ead2493d0b414b246567",
      x"dd7a2d48a1bba1a46de0486850f61e271fe2b27332a8f6b6d13e337b02280748",
      x"31da74de64ad096f7889a7a4e179d0863481d54f76cbae8915b63e110ecb2939",
      x"8e72380897fcefa9c849c1962413983ab08efb7058b1fb477317b69a4686a4c9",
      x"f4014b4c7fb3c628c43e9da7b9e043b134972f220cdedc135688ed874116667f",
      x"2237fa02e5e84d21fe17b83d1581d55f1f792ae91824685e313e1b46a621140d",
      x"f5d6dab21878c4b1b1bb6e2947fe0328de54f2d634629d58fd3ea5cccec6f9e2",
      x"9572514459b319d2c1ec50255a50fa7168cc08098e157d21e999bc4e99ab2e27",
      x"af4fd5b7d9a4e52818667855d86d1309b5163962185814d43b92d3f3ebe9d9d7",
      x"46dcfc3afa3b20d4caef0971d436b63d17fdf9f1e7610ef5b530eb3510243642",
      x"707fa0f97366a43dd0f4ce4df89ae77fcc639c8e7362480c9c36ad13cdbe830e",
      x"11aca634aa5e76f5ba37a00f7a068f69a20575b146026aabd39fcbfd5d0ddde7",
      x"a7f9d40d6441ab2a3f70dadfd9a43ff560901d622fe03d9f20ea0fc22110fbff",
      x"8e50744e7ac8be1cab6cf889d235fccb7dee9e8eb7e03b2830a3e9cc43e2f5ef",
      x"eeba1a707557266bd684667f21f30b38539b3f25ef93c7a0c7c770e52bb4db7b",
      x"33dbfc291579ed3ea7ee1253cfcb96cbf73d511117032444f56374941b2a19a3",
      x"802653ab0a10afc982e2f73026314a59ead5ba310aa52615e5fcd323d813e8ea",
      x"379d82cfb39850c4331967512e072cca6b8008d204dc3bb7ad5033ba8b1933fa",
      x"3326b59294e13f43917bfddc3e19d96d93ba04a9ffd1bc6fbee034ff346b2aca",
      x"3a76e194126886a02ddf968e9079d609d843ef9b94501aea19cbeb9f88addc2a",
      x"fcc65788a899c333d32ddd3e44a169ddbd6b2dc24424ad3c8b74414e36c004a5",
      x"e273a45869a074a16fbad071c72084f0431cc84d0987e9e493e87f9f89ebd4a3",
      x"b6db84c30d3eae7e26f3eac3e96966bdec1892905d8e8d502bdef97f81fad98a",
      x"0a34717a5c3d5f8bf456fd8862e30346a127045ce5212fc4bd1094ca1301f799",
      x"7b55e69ccdf17b7539409a315195c93a4b795778c3b1bf902e21dc03eec2d83d",
      x"3cc952e07e58a6777e8cce9c13555fcd073605f1ef8eae25d011c520810d7bbe",
      x"e23de4d469dd5db93ce2e9c616737731dcb85389d52af6915d29df59e8bee6ea",
      x"1f884610dfd567945944cb1cf5ba26f26a8d02548976ac65d233ff214ab637f5",
      x"1881429d0251f58a2c8d31f87f63225f5adcf2bd538474d7321b5f98ebdb7753",
      x"d3ca54d8560bcbdadfc69f6c7f45ad85ca9d73e22463586f540159e3588dec73",
      x"0cdd0946e9a4870798af8423c9eda7c01a158c6e69a6ab943c75f456739e31f0",
      x"ad902520e90731d82d04379997797457b142de1d89f0e4ac08a711eb7c6ebc3c",
      x"e1823ab42bad5b378d0897dc5596f63bc399c2db3b4efb805667f4f0c61a2cd5",
      x"0e8969a8a5c60baafa86f6ac3e22cc2086114537570a54d970a62ef1c4cd0bee",
      x"748c501948705d25b63b7643d57bc523cf86fcad830c13ce74340e5b4e30aeae",
      x"c6210c7b6e1d640d64b294f6e035cb495920287d1e89ac2c1afd81d75fe21eef",
      x"fb2a03b1b738ec05b9bcab1526d4ebe6142924d69a588fe2202f1f77b7699336",
      x"2a6d45b39e6e8e8600d9c5e756c58dfa1fefa68f0f9e9b2a9e14a191d315a670",
      x"918619c2f29c4861f5674915d9eb931ddb15342e2638ff16ca16fc6dd1960ea9",
      x"962fc1b621288eed493faca6a59c61cdcde7594fc0d6fa1e6a6a2329d932b2b8",
      x"a7f257da2e039e4234a684afded443bd72913083a0a49b081c941625087f6292",
      x"4307b61d081b3c070ea329ec9ad2cc2838190479a8cc7ee3c7cb8ae69e69c444",
      x"f554d9c9601ed841e650fedb96b98008c691c090f7cd8b46ff491334df99bd7e",
      x"cfc2d11112f5818626e7b876cf6e0c532c9dfef36795d0fc4f4dd2e357476b5a",
      x"e6998fe52906029dfe8ce2a12bea16059852b6f790f37eefeefb10298615f81b",
      x"7e4d81e87345992a6035092d9491ec773aa14fc7e126fe6c27243c356fc41690",
      x"a517fba1c2f1fcb2341efce5b3a10ba406fed0226eeea9edc3f2b93a113c05e4",
      x"b392146a971dae64a2cd40b2df38b6d5a646f254e3eef93700a4e243a6ea231a",
      x"5b744d74a2133a5129884b05176e538e072f1e2a7d00ff48fb61aa30b96c68aa",
      x"374fcda21898a9b694cfdac0cf76530896b3cb03a05fb1d6db1492a048e0a734",
      x"2ef36adf071add31c239087a08de7d2c5d014535348dc25dadbeaf488fc2917f",
      x"c493392fad6c48ec4e975e2b7be27d30354c3cab1591de125b86a9b048127e68",
      x"be64cee4ec91b432a9df384ad78c31cbf8799aa9b16e73e80116f6eb59088661",
      x"1223d40c04dc555adac5e76e19c50cfcec7e6cee20f3bc362bf5c8ea718560f5",
      x"97c33a49ebf35a8da889980e3b7edc4408a7ed1e886812e3ab3dce3ca66bb86a",
      x"0b46734884b0ba9756904c9181abf74dc4a985a19dee05410a2ebfe4e5bff626",
      x"19a5c396f89aeb9d25410cd90797b4cbfb88b95597d384945efa01325b4d2461",
      x"5cea08b9bd92c1d41afd4f133cbd9fda34a593cf8a3109c8bcaa0b837991f2e7",
      x"9bfafae492d6d2a55f51af52302f853cb54fd47d70c2a05f82bebe4750bd6e4b",
      x"d6975a75c0c465de0dfdb35a29cbb73384da603a20de75a723363f5a0e65118c",
      x"746b55d5e88a46d4d64336de010a713df04ccb193773dcae04453b63080c1170",
      x"a2c430750234406f3c7732af6fb16db1b4bd9c6c119156a06027f31ef87c2e08",
      x"8814a0e54db31a813862ec980ae4d0220e44232a494b7f704ac3ca1cbb7b9067",
      x"668d9b161091f8e20034561689cd0e0a7c5634e7d4ae0975d0a1830683af3f05",
      x"60f119b63c9d0ecf889537d3d3bc287c35e5776f414e30150bd9a98658a8a1b3",
      x"d5e911d745dcb401fedceb028c1209c8cef81e441c7b5bc7a4a440b5affbdfa0",
      x"dda9d85722c0c6825ac93b49bd71cc0fb2051b3bc7dd313f3a495a2772a1d9e7",
      x"e0f36e851be5fa88191958ec884bb150c279421cb36ca620dfa65d772d9fb9f0",
      x"60c4046c9002a1a274f2788e1959801b83d5f34b5e835ded182245d77c13fc00",
      x"da9edc0f56afd1b245b4fadc8df1611ad42effaa8cc6d4853295d14edfd10913",
      x"eb8e02b247b3e015466d16b8fefc214432974e57b29d69c0ad538c66a589edbc",
      x"1a0d9a6777497594e2f16cb1e685c1cf5605f2c9026e789904e7f9db081990a9",
      x"bd2e41fe9cb8bf128310f29887fac673d4224bcb86ff22fa77faa0973df18afd",
      x"20a2e6a535c31499d9899b75b469ce751abda95be65f75dcb474723dd4fc9d5c",
      x"1f5b3cf67f71ad12c3752615f8557c9960368bee67cd270c23f0ae62c6199527",
      x"c433f76115f0c9be72ea439544d7ce3cbfcf30e4df3735cf659c1bdf41917f16",
      x"5efc429720a6bade2ffb2c9275cd312d95f913eac2fe441ca5c5545717218b25",
      x"900570ec23fbf27cdc44ee19146ac6c26195ad2112fcf7dbd4f6d26ed5043f74",
      x"b23b8f6084aaabb8c85ac496b3a57c7fdfe75c75d661a67402385c647d285505",
      x"baf31e7a0b41d978f6d61e23a1ea28cf91b68a1e9f5c190aa6d407cb133fdaf1",
      x"900242e77cb60d99ffe7c3956dd4509a80ad2d94da7e5f53fb7bc53aa325c199",
      x"6cd68aa861189432605ee82aa753e9c9144930601c21b848e6593b9115923ac0",
      x"3b02dfc396f15039d389f43845f8c58e8158e881c1eec829861cb1abdf612084",
      x"016ca4c53d320102253f5097580ee0ae0f39a7bcbbb629fed6efc581aa01709b",
      x"b7286c106985bd7689b414c3375b246f7b01852935f699db19225c8a43a2d268",
      x"a93bca780511eaa4503f97ede18830bac5700386c518cceb4e4178e76d0cea29",
      x"7fa5f83498c73cef6941c91cb5c62a27be9679921abdcb0a8e6976bb82a892bb",
      x"79a6b666a94bd5c13ad5012519b7208e6ffe0e3ff78f53b6f61bab08e02917c0",
      x"a5430b700e3cf7b062e426ae4dea9741d9f723f1871743a5f7b17c17794687ff",
      x"8ba52c8ac90d0a78ce1201629c208a22733e3929ef28f2772be2feedf1ce692a",
      x"01ab710c0836305fc1b77cd23784615924737e6e5f1a83454ff5ac5808b0d6fa",
      x"2cebf2bc6ecda0198fbb885abb80e4cafc6361322d3fd248e022244563e96dd5",
      x"35a5fdfb28e0e3baf300123307d33071e1fdd9d53af041608e909080d4caba52",
      x"d72609eee24703280aea9d6bf136c8d2c0a48c1fa0629c78eaf98d53c5c8c620",
      x"217d855d5f83bb06993d75d51a06843f624fb61b526962b6ecf6a60d9d4d0fb6",
      x"6db3376048d9e371387511036b2a7f1bb6873893eec453b189d6ec0909a93f50",
      x"202eb78deeab934eef2852757caca95d591ee09233be231736536723e59a5104",
      x"b8d6f05c832cf248840954dcc7843d4090a565191b79f0097cedea60c3133bad",
      x"f77a33045f8511f59ee9d51e25f98217ac2f403aef54d282b085ce73b5b28b4e",
      x"2a66222d998c8a51d22c046237055c73b694d6fd4d8c7451eeb26379bdbdbe40",
      x"b7fb33f58ea57510c32c0b8b441c92c38d64db66fdf94f77ee622006b74222b4",
      x"a4288bc155536a0a307521299f3e3b701114450c5ddede45b407fa6379114fe1",
      x"1b6868901bbaee18967fc899c66fd2746296140719e3dc787473446a06324f33",
      x"ac85feb5418a83aed888a2c71de1ff29b7a29ddadf81846c6ecb26dddeadb97b",
      x"1f867dfa797b2f6db35c836a912d758e614902d2d3274adaf2b9720acfeca4bc",
      x"3acb7502144e487bd5f2f51de1c7336b86c8e8df00f9f44239a06ddfa0708f38",
      x"c3c77a8191dbb50f9348e25838c39e4a110b6a379ed979ead9d462ac88973ecb",
      x"df8d84745bb1b1f834c01f91fd77e52e8df89738d43a51472263987e6edde78a",
      x"d8c78d0cd97f316276bcc925f700edd76e397306e63ad5a05184d4d37c6ef99d",
      x"3f193d97bae979b96093f069da6c858749afccf7c859f2fc663a2baa22bf0100",
      x"cc816cf9be7db954b6d3d2d7c15407c1aeb8d0564b7055a47e728d37a6f2f2b2",
      x"372ff15f81083f366cbdaf52b34df961b28994ca3a90dd0d3c7ddfd67f92c931",
      x"5d3a07c79ac5cf8991670beea2d0d6b37c81bb9a7033ce7f1fb821625c207943",
      x"6e3cf5100e214d7d4022911cebd30acaedbed9d2474cc61e405534fbc233017a",
      x"c3db96c07f21d8c604b4d0d25510976f1a17eb0a47de60a3525d8372dcb58226",
      x"cdb9673816a8bfbe03d58bf6dd5569e4fe0399bbc050d139b7cf2c92355e4398",
      x"821dc36bc2f18d1389293bb6be7a5cc3af81e6351f71b6aba8349e08db5cafd5",
      x"3aae53d44fd1a12ad03b19d3d4f98cf8b3a9dec21415c1d901cf9d07aa862223",
      x"df28e18d683f461bd587fd9bce561fa86f58f36bbe968f2cce251582bbeb750f",
      x"0cf700e1e0cc56a538f8d8a693c84a0c1ed5582c16c57145c098cf7d370d3b14",
      x"cf22a7d0bd359fe9d21d38d2bf49f94488562b3cd4268bad96b6237a751e79bc",
      x"9e6cf5867f7780dcedcb05781f3dc17075f9325d30f109262bc5ee2715d4aceb",
      x"d8bb472d320c2643afbba70ef05e92e44e3758339e36bde099ba329ceda7b558",
      x"b2ac7bb85d7ce0afd61cedb5ae9ed3f51aa6fa52e92ff4fc2b4b4dc8a8f1f2a6",
      x"599ecee80d6f0bb95a4c7fc1257724680912377f9b8f20befe192e7cbe0e1758",
      x"7aa86d1d86a21af1418b759acf4564635f442f69996e5c2640b27fd2ba26a9fb",
      x"c629f5e3d3c96f387e6dfc010f2e01c2a38aadd775a02253c9dd02e7a0502872",
      x"3c3cb4461ecc972f0db04b32843ea2b0a234165dcab7ba9c8b1c3dc3fd1e7331",
      x"7076eab9006c8ca6d2650c462ee8403440d20633c80e82f20c6d122ae4915610",
      x"a226ccb692086f2a82b1d48109932516afac404155b4460efbd2ff155148b096",
      x"aed8a1ea659e90c3dbdcf6bdb5932c0178af10d8982dee0cc0a97c3ec981a345",
      x"bffce0c250b4fdf9580d966320d2379893286e420662f9588e9d8a1a033fa669",
      x"2e1906bff9c07a8b29631881b97f6fba17e5505560d86b9f88c82f9142f444c6",
      x"7589fbddb0e9f07ac4574b2b689c0edae8cad1d96a18118cd80e24c82ffd6362",
      x"2b6cdd91df69a198c96a790794172f0d1a5790627cc95a61be82406894be584f",
      x"f1242e563189336dc97e196ec041cfea1c966d2c4d33e5fb262f8ce78ad0c3a0",
      x"3c81c7c751e8765f2d08265975ae086e1809f20dbb2ca4a6e7ce483a5839cd43",
      x"109b39eacc9884fd0f0e5f5e722f00286d74d3b086caaa6ac3325fffa51dfd7e",
      x"9c1ecfa482691d9d5f86add597d1e42c0446bdc6e3c289fd945a8aa37bf129a2",
      x"b0baeb05c6ac31a100deb53e6e6dc289c0058fea537b2722442a962de5db3986",
      x"3b3214124a216cb43566fee33a525f79d2fe6dc061e27c7dcadd4b3c481b6155",
      x"6b47341ecbc116d19d2fa764024d586e85fd6a70f0872d7da4041cba8793ac5a",
      x"0a05b595cd7f6fb96aa80b8b4229a59e86f3c62fc9ecf3910200753898122259",
      x"11c23d3da1d340b8d1377e110c655681d9dd587a6a590e9000cf08e693c1e991",
      x"28fb7bcdeab573e862c3afef31b7b2a926ea807d8363bdb55ddcb6fc5a6f384b",
      x"d8a6acdd24ecfee15ebad0b4adf5853cd87533e79d45c59b629c3f3d0bd87d72",
      x"dbcbded7323b884ea6e01e1a95cdb7521ea1d028eb30e5087ac0f1176cef6f43",
      x"199274bc34736221bd1cc245bd054036bf03e79b51ccabe18eca36bff7d786cc",
      x"7edff90909f449cc082e895226420b13ea42da2588784ed305a96ede3af7bd4e",
      x"65c01e0bf705a419d84aeb4aa800e86bceb5bca7d8adbd4555cea9543a509340",
      x"1f044c4c2bb7f31edf3e93088ed2feba3b667279329ce18f3fc222c996dba419",
      x"d50d0d24b6538e6cf5a5ba0e7962f3d2aa13742d727b72373231be2bef36cb6f",
      x"e8db86765b1d6c055d91582ab8e7b53b12e9b7cbb0631fe81f7fa35511766552",
      x"bcc4b390c32057b13d6277128687405859b7d2596b0eecccc7de2d12c8865f84",
      x"49cbfaed22dc58535d31a94b471be84bac8e6490ea59dea85f827d42f71b101d",
      x"825c6c09b9e500c0481884c084d6756b69e3d769ad4731609de252e26e0219b8",
      x"c114dc60cdd6d15163b122d9970f7bd12dbbdea847f1ecb69b4f5c8f3c536779",
      x"1f14faabc9ee94a4b03740f5e1deaefae021920f7cc9a1c094d0b2006342d568",
      x"095b0407ec77cd8be0e29e8e331a6f0dbfd883ca905f5520953c12de69e77a5b",
      x"02e00968fb645b1d74fe97b9db192aca716f18e2af1d20eb910b78b599a20a3a",
      x"cb5a6a0e46948b38852b0538fc85f9ca25cac93204e0d8ffd6a345cb4125b351",
      x"b694f1af39254c9500e74386842fcfc42e95046661d752cdb1401e2aef3f37c3",
      x"d0da0da9ce53b19299dcb9f627c945f18cb2227929a9d69f394f4482e70b6f0b",
      x"0601cefc40e45b927909da575a95705da008f8b22a30c9f2cd62468686267093",
      x"aca1ff61b42697b908bb2a7f8b3d7d2b82ae5c13fa487d5c14cec94c50b114f6",
      x"829a8600c1a437ea82c1f62670469d2e3bc40e7fffaf3e467fa748ee8b1a22f8",
      x"e2c66b3a9ff4875f5310e9020ccc9f8f76ec60a928950d0a477500e404774eda",
      x"37b932c0d6bf6ac6c6c560e9834b01e4d0a5b7912b58d473a2cfb983b2647ca2",
      x"5b4496477d664a7f76723560ab1527e14d17e628f936ffaedd37f98e52ad9b37",
      x"d595e5e8b4c0826e4da281d55e60980a6b8da3f356d28f8dcd0edf5781fd48a9",
      x"1762a531f80f2b8a6d0917ac7d02b811410eb2d6746b06feb7927436d1d8175d",
      x"30ac97709267fdac8c01f946308538f8ed106d158272b0bd52e3153305164eca",
      x"042ba0e9a77ad1806654fad20d1eb46324f8cdc967536857383e4a5f0652877f"
    ),
    (
      x"3c73867b49478f6b584e49d546ebfe41e137484b82ac2da431eafef823ffed35",
      x"c03c33264d5f4d6d13a0e3fec0826eaae55b27baf38d19768c2bd3bb9cf0241a",
      x"4d28a0be13e9aa405d820a8e70de1a8471f360cf84b18fcd99130de864f703ab",
      x"3bd0f4edb381fd9db511b691b6d599ca72e666cd3265265fffbbb5ad724c14a7",
      x"80871b127c0496d775e4cde245cb513d5f13550549e6581d643ef7ed008794fe",
      x"baec1681ab5d2a3c3a296035447d0f71757bc00efbf65c97ad224cd37f22d3cc",
      x"5c561f7c291a94870b27dfc97538affc2a348d5d33c2d6487589631ab22b8417",
      x"d7562a441d27d7469dd2733f8c8b64954f67b88c49fe1ebb03b20e0854976b2b",
      x"09e52c1ad783f2e5916cf36fc1279c150a7e4eb03ef5e71d368910e1a70d11e4",
      x"e1caf64a67c14e2b35ca26a1998c6c329d5c52cf7cece13ec97e7ea52a39a632",
      x"e752b5652cd12dbf3673864b864fd4e922bffec84724aa21a4820b99c7ab3036",
      x"63e7d1e3c857ede36c79b4f0fc5d6d7e36dc47ae2558ff7b37f408c64c702a67",
      x"01732f51a4d63a98873eb16e2bef26b6848371932a96d6c3543d5cc648fc28b9",
      x"8946c1a04b15903e05ecc9dad1df4858bb3612c4e7cc9fe3f55b06b37d159949",
      x"cab52261b678c84e7d6b12a7293a59a9a8d2e5ea22001163fc2b9db0b9ad5421",
      x"cdde4914abc5694d372104e40cd69ece41372f4b407e9598eb228d2bed5eca61",
      x"194c3926d8c17ddadc7adda973b13f979f2d4170879718de9021ac28cdeb0ad1",
      x"e7bc1ea53ebfab88094c24e2369b0338eee8890a44b798ba96294b66643b63b1",
      x"1782edaf3fe139a59a364a82969d5c81039d21c2b860744b5551c692b38ecc23",
      x"7a20a7158acb7f1806d58dabacfcc50cc1a7d4eb6a77e11d5d191a170fa9d733",
      x"0d47cee333d2b0365cbfdc114f4cbaff0f6f134e619fe140b39d15719c438b73",
      x"a0732923bf07bd62e9d34585f21dabc766e48da4f6c4815a09e6bf50484f8b24",
      x"0b32cc3d261a632ba1ee11dbc00da2df01ce1a5809a406b37bc20f17d737ed00",
      x"033a1b3b78eac335b2d7b62ca53d194a6c94a3daa465fbe7dd937b695c5df326",
      x"5a11d4dd31b7d3655aad56dfd9d50b94991ed731a71c0e3110b1430ac590eaad",
      x"e665e7a99f994d4a2d94ae377036e9d5024760b055e672eee23cef5b74e0006a",
      x"46c8bf20fc6f0fdb4a2e8fbd8043c957ddc312bbee3cd191551ea2425c31479f",
      x"fc787bb0936118929140396e46e15cd23f017729893aa2fddaf043bf963d0fe4",
      x"6d7e9ff2fd2c2d0926420019d31d8c5b439875fc01ed2c22ebef11d4a6e6d7e3",
      x"ec67f2201c1e7b9b5bd65478088a3c1e5d8df593a46607c8d2cb3981c9f960bc",
      x"2192e66bd13f8f7d8cd7064639de066bb696d673a9fb0038b4b34eb88894e2d1",
      x"ddda3822a9de0341060f14c7c390f292ea8f085c194ba036d885cbf01bf4c99e",
      x"f0d69cd1e1bc8e5128177af5ffdfe04f968afceb3f9ee98d072d8173ab2ee8a6",
      x"b76c9646b40adeb00d96070464d2bdba21d906716ef6fd974ec3a4e1cbf9875a",
      x"e7b7852b9ba998f35dc2a59ab2682192502d76f12d2688d833ceb95bb5421fbc",
      x"2dd6d9bf462aee7206e1cfdde72aa96ed2e9d7dee13992c30c6294fca71a8461",
      x"b5f06602c32dcf92353e217e7b587685e78344805d6491ecda4d61b7020793fe",
      x"9ddd68d50abceba044faf8bb7826406665212d6fc0972e76164fc29343e28355",
      x"89457880db10df40a1749f755dca0839938da4ea36438531a8d38644f53689cc",
      x"064a06dcaaf784fc41f1f6e8713ef1f02f6dd7e8b59b7209713590c0058aca86",
      x"06c50423ee3db617a280f03701618963461e211603bb639f96c266341ba68b46",
      x"3391c41352c51c0270fff4e0eb1d676a8aafd6681bee5c6ff771fcc1d8be361b",
      x"942658f95ac794362a6286d3bd23e58977cb245defbb9ae97ac72ac7ad895e62",
      x"64cbffda9247311b2a8773cdbe4358ef09f54e125b3cb9ab50cf14ffc4fd7dee",
      x"2c973b1cb3ba2d9390de91a89baa35aa47fd37356391c68e225a0457af218de1",
      x"1ca03aaa24419c1db692b7d27a424c86755b290526a28f1bc76a3f87b0c8da79",
      x"8d68874e6fd6e6239988d1ed93c78978da5af96afd62f964e4496f30d41b4745",
      x"7640c2068776457c3fc41645e9f9da6a0a907ed477a70aca749e914ab5b5bb2f",
      x"8112d8d4ba727b7d54c7f163a597e51a658b0719fa092c399e202eecdb50fc2a",
      x"e29c6b14845b4bd3bf9cc0c54062ede5ec98722f2522f8ff5181541e10f2ba48",
      x"761182d821f239aa8710468acc5b2d56d30d05b7b4784d6fd3d9079df041276b",
      x"af93cdc44cfd6c5e52c74f06da7eddcb23eec208b1a26c18c18048c97a480965",
      x"f93872db9fab42af09ae08848cac7d3e9fd73638208a2749d75e7b51195a295a",
      x"7324baf88df17ccb67f1a89253bc29e5dfd4f85f10387938ff4c8af661145838",
      x"e786955fdbec3ef6ce82bcc3067625222871fbace5d47771b216db2c1b8bb31c",
      x"a4ebd848c79e1bf0f9c86df1c8777597ee0f0ac91ee280a12f9966390960ddaa",
      x"2ed5ee75b73be6b6a2bcbc3b33c8c4f38d21fa2687eb446fde8f285be2925b60",
      x"06e1863ac3082d3909637c91bbde8520a450b2d89c1af4d40955023ffca3d941",
      x"0081f023dc8c8e72b4e4e76e092c040046f5108602e7bf3d39595c915bc9b04b",
      x"d2b1ce5a084d200f867d8cf63c8ab75640c7a450643af252241e01d9e812f891",
      x"2255758571c4b5648a4b19813ad7a4c42a38fa9541e36d35e03eb32cba1c7c28",
      x"87400f48f2d81eda37c66093a6deb7ab2e44b51f99923cd59ce52cbbdb4896b3",
      x"334a9f392bc237441b10081ed72fc219559ac68cd25e5c296769aae25b96c40c",
      x"04770f08a13310cbf2fd39324e3c742de2cb3c0f4c60d3988544f054df67f3a4",
      x"6074142fe85f9b295f9a5005f8a92761ee1eaa22dcd7f546e2743dda650114e6",
      x"307e7b85d69b692f3adb81ab154f4b642818a17c1340fcb608c988ae2e6b4f63",
      x"f1a346ed0e6ef07871f9a4ab410ccc5861f87c7ae183e8433b6c0f33fbdc2449",
      x"96bcb6da8fd2e43c1966346744454263859002b60a1ce8cbd8b83f82cf5b548a",
      x"15910cb2cff6d89a868f33472e6af3e8566c1fb7b93142421a4f22bf995c2b33",
      x"5e7188f7d93266b03c68f62d970a06a4a0c653eb2d73ee7b4bb85464dbf56d62",
      x"5c13ed02d017a8788d2c1e7406d8bd5e77bc1a61a1b42a813ed7e80b2cadc87f",
      x"4f35d9dfc4845ca2ab7e5d73e821dcd0eef7b3c990932d0d22d2d224743f8ff0",
      x"15826652970d22941da3cd0ee7c653a64ff5afed9a17c06527ba689bae7ab035",
      x"01ee5d0825ec02c8e99c449c76dcb3fb21ba3c16149b733993a5ab1231819c7e",
      x"a5d930b58374c6d43b2a1545731649a6f3e2ba9730d734f47b42a7eaee0d8a4b",
      x"eee4e31ddc6995ee7b3e99d95ec727db320e96fc9f282feccb5150b4a3cd85d7",
      x"3b83dc34de6b589661721e882c71f4a4e9b3bd59e5ac3c83d36e9da3fa514c96",
      x"9398601e6cea6228a73bd779ae0794078d3cd5db29ec9513bcd904bc55b3a7b6",
      x"d608f49005fc405c5384044091b43231938eef994589745f3b4951ffd2b0d44a",
      x"660ba6622fea30fe5f2b47a0c7883c8f9a3f1f7f418ba79372d1080b3d40c21b",
      x"85072b4477c48595f57b6836860ef1821f6921d05bd546c90d18dae5eb7b6bfa",
      x"a3535e921570016a50ecbd904f0ebee9b272a5697307b5976012c171d5f9d661",
      x"f054b9197df997b96b42913c37c3626ee4e9190b68a63d1cdf735b52a714308d",
      x"455e73b95945f93849098d4a4a62e00f7fbc621e6f242aa533f835b5c50f26cc",
      x"740162820695dee89e4be2b06a2be4cad0d2888fb9b5d178600cf2b4e61a047b",
      x"cacb2608b838f1efc49b99c8023ba6643fd3aa81766a1541453863d31bcd1177",
      x"243173394f02042d6a67e792a90ca485bd9679a193c9a64b069f3eaba9920e10",
      x"a23de56d18bde757c86e6403c76665edeb326018031fe716c543ad701d67855f",
      x"c636e9d7541508aa51bfc0bdf27877d0a3e295356413f4a4717d3ac4fe9ba5e0",
      x"a9de45c353676bf154398551031b669e0e5fed64d8dfc699d6742c4a5b188b61",
      x"47f4497782782fd0c725dbf928378588225a96aff97a6543a65e47b0874b805c",
      x"538d34369603900d5073983b133515997ea4df9b46a3cb19b03babd5d2c354b4",
      x"58377a1c7d6ba7705149d9dbd5970471ae9d0fc7a4665705fca5a79838bb1a0a",
      x"7e6c207dce9420b641cefd57e8b6d8adef55ac70ee9d6d24c2f085a701db76bd",
      x"aedc12bcb31ca9c0b93bc3dcb5098fcc175f1b0ac0f031ba3180acd2c594457b",
      x"01504eb310c7eb3b0f230ffa5422817fe798886ac288fa9175bc74b651df3e29",
      x"6fb68a6396a71f34bbd96c2d4826bd6d8beeec12d5a93af1c217965043f49f05",
      x"0bfa6053df9c0b00b01bec40ce7989184a733a52868d22b703dd74275401155e",
      x"d863f71851b66b8a518cdace31c7de1e7fae71470c809d3dff29b9da365b4911",
      x"8939e2bf6218f1e82f76af76a7036093d4a1a1b0734b04527339112c33196172",
      x"f42e3624f5cc58f6350d936513692396ff68c6eb9f0a45737ba0a492b28763f1",
      x"d6799c2a5f2a1b20930ce74c32782f3e8620e4e859cac1f8a217e8f2df6c64b7",
      x"d02fd17d48c3563c62952991a738ee1434512da93a65fb84aa0ed7fb9733fc66",
      x"a3861b85a28b52c1a6681bddce1b3ca6086202c3f6d7f93ac5cc5b263e3b2dcf",
      x"02ecbf9764b351db68e613405de04156098fb2029f843cc7c0dd7cda803de5af",
      x"03ea91f07bd28227511be9432095b4c0305b92bd8ccca932b363f8f3f7d1e1b4",
      x"84ac46a000a68e1d9a3f93a69cf75ada0c6416fabb332f4eff647990f6f1b898",
      x"9de7100b15dfbfad22ef4afe266a95b2215fb03782978a5b033b99875f796e20",
      x"da308d005026d047be2cc94d876a8ba7a527688cdaed2ce2c2a23c78e977bdc3",
      x"1e0f661ac53cc3e6ad02ef22dd6727026161fe2941ed5d22917a7ad5b3668b3f",
      x"e90253f98e33b737b3f1e1ba000b88f6188dc8ce990b721333dc21314d67f86b",
      x"4d7e546d30ee9f1248596e71f7233eed553c3cb795af7e89aab397e4830f6055",
      x"19d1e5d3b275a73de794ee91b67bea37542969163131d96aadbae9ed4447044b",
      x"604ec99f2019b8f6cdf329ec7e98fa8f6c5df9b65aea1523beb1dbe571e9df44",
      x"ac018818cb1a1cc9391708e3bd8eedd8a8f76f8dc3b8a798398c9481444196bf",
      x"f89a94949c7fb8b39c498ab4d1849cf12a5c0d04cef622dd2f3eedb8de14bb9d",
      x"fff3e15abf40d20dd45fc1da3bdfc38806759d2b72000b5e484360502eff6bb0",
      x"8f6093dd982f20d1f724b4d865ed1b5e095968491097d264475e951da72102f2",
      x"c211b8789a9d2ed012f29e7a50c01c2e76701e335756323b5ca57658821e761a",
      x"26f374b4d5189c8c8a0a92801c858ff384a774b2e84276aebfee1ce89ea2c681",
      x"cb5e444c5a1d679a8210227684f41ea680acc47f31dfaa1693b27f5267551e0d",
      x"bb63b2484a3935b402b1dc5662ad6b32755d5d3c0537e1ca2cc7a4b760bc4c23",
      x"5d43a7212243e0f572b955d138b31aad63c3267c96eae6b1b072c837f37ce493",
      x"46958964e5fab2febceee909e9c2884151ad621fc2841526e1198f6df846e8ae",
      x"2cb0cc738d4f646e25b5af13c6954b5080dc771a29d04a0fc84c941038bd1376",
      x"6bbbce00fcb694badcfcf4bb982406b4f88f73fe980896c1df4b5f388e1a21a0",
      x"b7db82478d6ae98556bb423f577f7299667dcc1960b53d35c8d030b6083d481d",
      x"5418538ff8b9d1e0776c3c0104343f1bd05181cd55032fe6b6c4145ad8669021",
      x"b69cb5fc547b1be4f3ff7424b26be32ef30ea58da274da0f8858d6f47448e16a",
      x"5de0132c43ca18a25e28020d94a4d37c6d4ab41f06cfc129aae3c2397a5cc116",
      x"cacb13d79169a6684814fba0d81d939a1dd4701e25683cb5db239beba198ef98",
      x"2da271d28af0e0e352a6c4d495e54dfe658e22d9502fde6e9f1b27fc25d49148",
      x"dd9b809817e8020c5ed4c332f0b521a8e4ae5ed505d4808db7003b213d69af11",
      x"01c0c68991e10e00bc47b0e43a9613fab05cc8756d45a1af64528f05e7553787",
      x"f0047e098269134109defcefe5fa1a33a9114e883b4277fc531f96d9e5ecbffb",
      x"c1eccfa94ec81dce0dbef0c081b4f65074d68599f91d4c6eb204c6f4c89a016e",
      x"8c41dc3ea008cfc501efce47c7d2f51343f868ab95ddc8e50c86573e5042a4b1",
      x"b81604bdc3792d765b3b3e762b4f834bbc1abe2c8f0befddd29d70e1b67eb577",
      x"ff27d41295c77a93276a5e5b97a364629db5e62f4e249dac3791e3bd076e3b7b",
      x"f6e702078ae3014b730eb0fb98090e9377968e79dff04a28e0539206397acd74",
      x"ed7d42235c94817359c03e71acf9c3ee79254e40d1c3f77083ffbef675528603",
      x"796a6482b3df1effdd56148ef73ca91c6006b80f55e65a10402192ad259fc237",
      x"03bcf148a43e29a912f9cd70477fe7e9f0157c2bbefe08d27589671ebdf905f7",
      x"93758097c2af87efb0d3d5a52dffea21066e9bee195628b54eadd319aa6b1be1",
      x"2d5cf6e3692e45c94ff845901b5e73ed410f6c0ad882166f370f76b5d109ffc5",
      x"ffe744f8d02d9cbad22635278a76cca690b2569a262ad25ff1bccb08489d36d4",
      x"822958d9a04b67b17ed07d05d3ba928e0e090b632fba30bab2e9dbc00be93994",
      x"a2ca9021a8c4c172471c0db145d0f4078c98fbe24bfe73c94e2a037178403e0c",
      x"80ba3988fd6cfb53a69a54771bd2d85f2f55836b221e0553eb1cf3d37c355a52",
      x"38642116293b996084f644c4dd1d2bf97484e537ab9e3b9981e52a925c4c3f96",
      x"1c381a6ac3bb0ab3e9c81fb9af8701452021fb2972ca57233d3396050a859686",
      x"82fb5210d51db49a8a50549fd2950794762559c621c05cc2e4f44dca0e5eaefc",
      x"a1832372fd086a70555b337c9f62244da47bd79b9b7603ddfa66380dc18f6936",
      x"e645bd7f012ad6f8f6afb5a314327ac1ef42ebef38b4b651226287a784b7a444",
      x"0535e75c24b19e34a0b7a1f3e5c1b04e07b017beb34203b6bfa40a8c134d54e8",
      x"45ea5767da86c89fc96c8797c68a9b13fa7e7b68c145b3ad4ecf3d970cabd6a1",
      x"3e733b1b853046461ce44460ddbf247e0729b05aa6a50fe553c9d0236b71eedf",
      x"df62cd114ef12743b13424ae0ed506682e4cfb3eb95003e5475c8b9fc0d58aac",
      x"e824df81a01481a8465c6d2a48aa41f295b32fab3b966f529e461e5070cb778b",
      x"097b5919f5fdc2ad7e7750274b05969e8f52d9672d7c1d2208cf2e0ddaf1fabf",
      x"fa9d725fba09543e1d753a4cfa0fd005d5b71c063131fdedcbf318720663e653",
      x"2b5567a21eff197e069f591aba917c159bf5ee533782f8e6e01a022eca698c81",
      x"2df693d16ea368e24b1200e061943cfcfdd9d737d10a4155ac85f54b48533724",
      x"9b37070e8bf6cdb7930d13c075165efe8f53a00eb88e5d0cd658b62e20234222",
      x"0b409a89f7e970e6c5fcc2cdb461b6e0c1b930f1914de5ac785976f44fc8ba59",
      x"19ca3e0c53c9d23aa4e4db55d343f2d95311ce10c3155745f7646f6fd0b3a1f1",
      x"840d9e3e5749474d61bc6a648a5f7aac9b397a57f2503cd59f4c631b59e0ddd3",
      x"c762c628593675eb885c6ad98cc5fec37ab9a230c4edbb55651d5073c27abedd",
      x"1f8d3b028d7f5e4ff8a606df28b84730501aeb40276d57a47db3afc824ac80a1",
      x"5536dcfed08d694794e8d34aa9eff59ff1e5dddcecd0fa1863b8d5e6a4f40590",
      x"88bbf6254933a26d8233e2ddc367bfa39d44d459ed67d7248c13de7968f0b530",
      x"a42db790eebc6f54d21d66f581933e21d770633d15b270fc768f6e979b2d1157",
      x"973dde6669ac2c03bfa73b7a9fc9d83940c197d4bccfadd173e7869946641d69",
      x"5e3c3d3a895c3d9d418319785c3d9e0de7a35e7dd48d4c7374dc9fc80f1a612f",
      x"f3ed4b1bf0ac70e100b3c7f247c2b8551201140156117b0747f3dfa45fa199df",
      x"2d25b5fa4c91c2623e6382b0cd2152358f29cc16eb9f67495bed375a8efb8717",
      x"55021644f1cfbf81616a42c922c18da57b68c56305feca919c49844f27dbc503",
      x"51be9d8f54c8828c780fcdcdd239656605a205fe86753b4a7656d3074bda66bc",
      x"f75950a54968dbc303863d9124544c1023e1aed6151a47a00d21830610448310",
      x"575b34af0ca75f15318770e7a203dbd9f18b7f8e231056eefd7c7d246dc8033a",
      x"a61e70987564ed98062c3941c3b58cafd7b6fc6900df488a802692c89290721a",
      x"00177a5ed1053c519c8783f3f303215f4768d5e53b701e985b2faa09c76c496a",
      x"eda9ef459ba6350d02ba1c2e8fe403f52da3c2cb30b0a6e14d27a5dd5659e8aa",
      x"c7cf8f038ebb9b62e03ae5c1fddc2fa316422cdaafc3c4ff65c96cdac834b22e",
      x"e9e1106b0b4899614bb3da2d9109752e16554c62d0307cc5020cffa5a0514e4e",
      x"c06ea039a6340b61ce980eabcda1979691592d34614dbe870ccb8843c588c8bb",
      x"2867bf4fd65ff0e175d356de3cb7fde1ab2006f30545cb35dffc35f15a92bd20",
      x"fae04610c3b009e02bcc99326180f0f11d5e0292d39da0a272882a91e4fc712d",
      x"1e8b6b30720ed8029c425f9cf1ca39ccf8ef782cac88ba38d319599665fa666f",
      x"f9cebc6dcb04ae885c3d3b1f4e28e0daac36a5ababdd1912a135507cdf29bbd1",
      x"4f6ae54475607573975d1415b7db828cddc66ae847547862cc509f41af099d00",
      x"5df7ca17dde6725add3cca18a892288715b2a5a550e220a7bbfab89a5392fc9c",
      x"0255c5d95a562d59129ded2f2a0b8406b0f2cd41e20d466928eca1f2e0ccd9a4",
      x"3cedac2ceadb6b0dc3951a96ba2f501679948b5c3d4e8927db5303f04bbc9eef",
      x"128a02a8637bdac4d8340fbb0c0924b9371a7833ab724230545ee63f63ee1cf2",
      x"97655b689657c8e8ff614b3e63d6822c2d9a3487762a11e0fd9eb07313a814fc",
      x"ffd7bd07cf4fe50d4dbba5b12478394dc838d994d29f2f421805e2b05897a14a",
      x"0136cbba212d8c2e57577b324812342373187ea179da9dc237818b838856f59a",
      x"ffc8eaa133ba8499b94dc4502afb6f837c72e123d0967af7e38af8bbe45012e2",
      x"d6d379fe859aa30a93686b5b2c97fe799c91afdd0e0127eb179a932780029338",
      x"0257fdeff928648b89cfca1233b18355bdc384260a0ea9e8a18949d642d45871",
      x"475198534e30b73b095dcc29635770ecdd00714229576891cafe99bcf2d54d85",
      x"b5f976bd71661bd7dd72b4d8a2f7dfdca47894a18932fc7c61133c0806ce830f",
      x"11e026719c95e871f60dc1657088f1299d20bcf7d6d94f3eca8ee8983013caa1",
      x"56dc7f0a86a5eb43056edc0de3d16e5e426bf0268ff7e719b3368eb1be795b30",
      x"3c5be9ee084dc5b98f63847162f2c3dc5c8696e305c533bb96d2d6e694010d43",
      x"226e43fe70be846c9807b6531ba7c0bb401c11d517175446e0c36ec04b2204d3",
      x"be5395d5713fb530e7ebd2d8a2a8071f14f83ddb04759825bac29828c8ac6996",
      x"030051fb68b922a6aa1069a76a2ab3748679bc6e5d6578ebba9e5ac62541a3c2",
      x"18bebac07a53538f2c28283f3863a0c356b45e7593f70d7c45c3708d1eacaf22",
      x"3fc3a06770a86918be1cb1d2e5e7cc94b72cedc23a8b42bdd85db53afc45e9f1",
      x"c0c4a59b79f05f29fcb9472593cad6560e8384d657cd03a8cd892e68048282ff",
      x"46ed5c42e8fd6e8d1c615bd5cbb632a5cda7460f1ec4db7a0ac4f4fa1b9a8ee4",
      x"3440488fcca82d01933ca09fc9f5bfd955f27b6808800b92fdcc6a5b9c0ad909",
      x"45ff8e2c7abc96aa3214a3f1a8c769c91add4c0d254b7447139513c03280ba6c",
      x"5d00c7e1af027ca15f80e67d503948a41bec3a3acd15f8f189ff95e35b93ffb4",
      x"034778be2dc48e70d612404d757531950b173e1ec333c949138ebd6f6824078a",
      x"c4c4ed805ccf49b62d0605a969e08b33e5eb6518303e8c4b2897e59b48c345b4",
      x"1038240fc1b8b0e4b188864fc52e50b3c6b98963207a47d908128d5e1054c1f0",
      x"3f7992a5660ff2505490798dbaa955318e34cf02de6d0872113c18444d7e914d",
      x"20f877af1622cb36571aea65a5e79b8742aa9641b58b0f3455db0763cbba4c02",
      x"81e7cdfed32dd98ab0c4fcff17c66c6db96fc3916f0c5259e611f879b364317c",
      x"9f06c073ee3a68e7bd3faad751b4e9ed91ac172f8bd6fe47c19b32db25fe0024",
      x"35fbac4833eebf5b9194505b03833cc349338f6de9ae85067fc68af7cd6b27e1",
      x"708e5dcf5702b15bd0c5b63ff81b95774b9352a1a39d59099513aac8094e8b33",
      x"6280652a405b57c28430c67e4cd889bf9160ad1e6ec0ba1f9f4ab7a755689c4a",
      x"85097b38566ea6b184bd5ab6dae805c2eb8d7ed1ddc385beea0673463dd5448a",
      x"a01d931fc656bcd2b5d54cfc7ba82b1a734436ad409ea7b68f4edf4aca3e6f8e",
      x"02055b3d06fc8d549433000d00e0ea4c6e2e458c490dbcb82dea50f365bca5c4",
      x"4931094f95f6312d13f4561dce556292c4893283ceb645163555f9e13f6f2abe",
      x"5678bd650fcf4901a7a7a3028b9fb5b6b63437f569776bd83c16dec86e3b4549",
      x"067d8409520c4e444bd6a375333f7b24cbdf9f64a378799d4ec38446370e4509",
      x"fa8d9a8d1f7f05fd75876eea47705730b754e9f7c75ea1367b68679115b9a5be",
      x"3eb3be50c9b7307803b297b74191547ef87a36321c68cd0968d5be00b22c9afd",
      x"5fe8b478c770fedd60ebe322b0d3f25bd4aeaa3932294e90f17b717aa11721c9",
      x"a6f3dd5fe74084db5ec04b67566c5ff8be534e7c8e2db07b7be06fc113bdb596",
      x"953d5edddefdd9d47bd652076b98e8f11d146de0bf4dc298b8e9d028edac7e20",
      x"71adabd50eab7062a3dba38578e98ac721a5a20246d11c01735a88902e0f8978",
      x"c3aca96bdde8fcd9a7c9c332cc23177496ef810b3341cefeebbffae1683d2622",
      x"04feb9b5873c7b751a454d2f97b197eaf1023125a1be7dd3c4b4af2805f58231",
      x"3e5f26610948f2f2e3a6af236d7752fc9a0237546a76d71c38457bc0576db6e1",
      x"8e5572b8fc4504a7c8b66487b2574065fd3389a6c3078aa1e853f8fe33ed8205",
      x"5da6206fb9bd8eb2e23baa383496d06b3608d7df9902c9bc99668a48bf9df1d7",
      x"132fb854bd96cc9cf991147a87786bd151d92f32f283cbe2739663f0250086d6",
      x"08ae214f3061ea33120ed46ac0903c78d0bb698e0094ff300a1459fd9bda8214",
      x"0d3a798126050129e60d6c25665dab0b504c79add02116225893bb5276ee48e3",
      x"5b5a340e672ecd429ef0f0b657de7d32c53bf42aa615bdbf9dccfdb0136e1cd3",
      x"772ffe96add9a9df309a2b4c8dc38a16ef25ffec89c5293a9d6e6d01f19eac6c",
      x"9d5ad4988bba724ff2634c0f52d4e7c72cdaeb6744ffd163865eb14ca5a6c2e5",
      x"cd1163d0cba6273562499475e60d2782c1b14084a33479fb29c934fa65bcb265",
      x"6d57e331f58d23af68fef4f51f631387e66f924d9d8dde5df43ffc11917635c6",
      x"3c4cd7415ae9aeb00138c56fc4f8e54dd5a587ea2984b370a290d781055be688",
      x"1d6123285aafd701c5e48370759ae9c39e8c751ed3f94bbc2d91b816d7248afe",
      x"d2d35af91efe1669b1c4ff155705269dab482b3c35fbf68e73727211aaea1885",
      x"d2898744943ec72566c827742bb707877e830b98faaf28087d86ae0e928c5f27",
      x"ebde62e368ca07dc5160498bff2596b2e93b067b0ce090c061b0134fc390197f"
    ),
    (
      x"138a3824a22766099954dfa4fb1fca66bda58911e3e58d49d068de580eb50ad1",
      x"723b7e186a8170f544425eb571ccfeb7db1fa1b50b64686612839124c376e02f",
      x"84757993fb9440821db4d0e456d1a0b4e3c65b05afd2af0009ab38e314d3a463",
      x"f2ad8ed9b733545d794044fe2127b1057b4fca98f2f3933d772c28c9fbc4f88a",
      x"a79d3a5fc241447b00e8a5cb1b480391000c77fd48dd039daf7283d1bdf5425d",
      x"260f89aef4343ccce9c8f8f6fcf13f9eeb57c76228c713f3f723e0712408015d",
      x"307058d2053a9c55dfbe591ee272f78cd2dc38748b0748561b336e0c6a6acfb9",
      x"5733b4693f058e50f2c4a92cf73106aaf626b130be48b704e38ee89032e48866",
      x"2ad5d78035a1d95b23c98210c63efd14edf2f292f4e6a64b41dd4b23073e5803",
      x"091b42758457f3960f827a415984293b5f66e4f60538a03b05c6f0588c636904",
      x"fac2c647df602c9cd4c1473712afc16a514d071fecdffe089a31176f5dac497f",
      x"d51eefd34decb140c85308f0980af5c790e8e589b17e3a4f17cb01941721076c",
      x"e28e73a17cfc777b489852f562884deb03b43c00a8bbeeefc91505b1a04daf2f",
      x"9c271bfe78a3c554d82aa6955e6ca44b8febb2b8d94412a47bc41fd2ab18a1f6",
      x"dfc1b556de88ef5731a8a72d8304f66d8684f311766faf7bfc491aff4c1a39b2",
      x"bd1068d109809182031a2af5044097d6c43dc1ef44fb11cc4b0eb1d257db6d68",
      x"af7d5242dd9f62a7791442af152b0a4ef630eee770d40913add06e96cbaf5d93",
      x"7e96193e080eb8aacc6e25201823654ef1f0c599fbe095c43f2cc58e477a9a83",
      x"0879a475a00cdb6a545310e6ff27247aef52e953098c3785d80a1935f9041d88",
      x"22cf807e2bf0474aa9f81ea37dd076f3e64c6f7b67cf12b5f128cb61af199d86",
      x"4c6eb19de8aa144f192ae52a26350715f3ba1cb7976b07ef0059945e1193b320",
      x"c903425c655884c54cb7166bea33ed1c9e0c8e3111f9f6d1ee09288569e47f1c",
      x"23a344a5e9be5e842d7aa03e26789d8c7bdca5eba9c505d033360199b47c53cd",
      x"5fd2004e79a58744edfe56b0e8f4dffbc9f710c19ec0d68be412ae306301a60e",
      x"555d5b3eaadde2ce1ac0ca4a5b2104fd9c6dc1a906e13e4285a4b5c3b5184b56",
      x"99ff85a5b599fcdca49d1ca6088e61a1e3d227f5ac9505b55d458078fd4f800a",
      x"b992bade32f5e44efdf65310187b09b86a14ce9bb7ee0076d353c7d8f4ebabeb",
      x"7aeb0c2b95b129fb34e881762146f763b2ec1bc555a3a13c2ff5d73653f7677f",
      x"728bef1570f8c3e9bd65342067a5df6f1f99de349e0c572d4e7595f0eededb76",
      x"c2e0762dce7ad281e5a1f1d8fd95aa15eeadb5eb184ca66a7f51cd153b9755cd",
      x"78b524a72879eb3fbca1e99257aef6d2f0d4c7f7065e73d04e65bd296134ec81",
      x"02a3d635044a67e9a229bafe20bf4a6a24c6e83b3c8a8f5bbbaf74388fb2ad21",
      x"197b2b68cc9f9f2ea6c340cd4cee669a51d7e00622ee88dbe2849f010248cf06",
      x"0ed796d81789af241293786da02465dc283467e25812ccfd216ae50784bb37bd",
      x"1d55ff85a2b7cd29ffa0882c0cd992b6e1c0e576050963760c0ffddd25867b0f",
      x"d05a3fe7677eece7e61d80061f2048d29e2cc422ad73f3411b14183cd6e43558",
      x"82598d186a56a8756c6be04b62fc01524f6ac6e3f752f6e2c4b38c4a961f4b04",
      x"e30fc6631b47120a9f5612ba45ffb94ae6d4d1f81a4394c20924f339735e8dc2",
      x"4c65b33065d4bd049de45b5bbe985d616688c0717600b2d155d7e2ae355baf43",
      x"6f29b458bc448410e8b1c5732c9a6808a3900f257bd69fa03e9b42b936a87e80",
      x"3f8291021c1406eb729c69ebacd6306578fb5af88c34e37cf3aedd3068e7c439",
      x"e8320aca73f21372d4cb98ba4fa4ea1247696c8440a8c166f1a4c3a5fe4a9d99",
      x"9157cf8ebc762c2ec76777f81e81da6245604931ec88a27d85da60b3b855ad1c",
      x"57417b5a9f9b90cb27a9f0336f14a993903dc82103b71084e4a5d3bd4ac115a2",
      x"5f4ed50685a8870abdc9a0193d45f7670b892136c4fe6cd74789f4207fff55d6",
      x"68ff1d1f06f8b50d2f849e4836cfb5a7f1b7d28e5a20a4d4df9262c956b76fcc",
      x"4ab51027809f3448e8701bc2bc8298b144a64f3e1d5f0be07482525c48919fe6",
      x"543d90033eef8d656ef1f2b73e91592c5029cb3b4d2a21cd65af000e7e73692c",
      x"cf03e1783b8c2747aa9c9cb462ffa1d9d5eb57410f781110bd1aad72c3ab9b94",
      x"5652788c54718bab7a76be12acf058237608f1be934642088efb036a635f1e23",
      x"872b48d92ac6785872ae2d1039986b1090d12b2ed1a14bf1b544dd666ac255cf",
      x"3186dfc3562189908c5c6b9469dfb796008e7b085af44bac5e6d6aef1145e87c",
      x"dc6e08d9d06488328eeeddf1f6881c2a39808dc4e91fd3c9fa617857983a6c2b",
      x"9cf69690655e3516a6ae71204e10659ad9f95aaaf40696b696ca47cd4cdbda10",
      x"68b6898f45293dc410a235e92b0f719b487d5895c5561f51ba33ee93d363c814",
      x"3df3f9f68b03fe9ac4310cdb098b8fa52554c741642e58d9534337dd74a7c500",
      x"b2b76e7c053b77703a03f0a66293c6451f50f338db984758a2df375a14123534",
      x"fe6251cae7b571874b637da924f96ef94f2108097c3e0a7d280ca9c066784996",
      x"b0d88d91a8e61ffc3844c9b9b4d6d01334747cc2a35e90d5a5d9c30bfb02c376",
      x"1c48fd8ad9bf5745f62fdfa57a7e9c974832c29e4c1979b73b4ad31ca17cf61b",
      x"68b631bf92f974677a66d22a5d4544c4d6504b8ec5bbf63ce227de7427b38bc7",
      x"a692daf630f74bac52e6c7eb96f3f101b0d176e8282b024187660c4a9882f897",
      x"f8f72ea712a595a35632ed7ee1e3509a30a7c9ab749ac9bb8654c6a9df52b17f",
      x"c85ccefc84518d97d26076e5e93999ed1f5d7c479fe544f829947fc8d6fab560",
      x"c9d5a04b6723c553639bc6263b82e370f0f21b507cbc39c3bc2bd545997e3c19",
      x"f846b429e4558eaf90853d0a90e63fd22d7b37978613a683caa4a33a875e1fc7",
      x"a6015b8c5aaaec8586207080d9c1271a4aa5166df3166f768ba4022abed6fe31",
      x"7c700957f2222befdbdb6e97ae7f047c4e36711f0cdfe2d6f4c48c72133fca34",
      x"ceec9aa6d2aeb58c75a5da761c3475ed3c49454bbe75cee3653c78482636c8f1",
      x"e97373d290f2d5065550af7dc64999f5c080bae68db977595d0a5c6dcdcc0365",
      x"d065b7eb2d6050e7d0073c7133408322212fc5929bb5bf07335e200704268c32",
      x"9dbaaae6cc37b998a0346419a315bbee43acaae671a94db8b191c7bf27fad105",
      x"b37571bf11b32ff79fcd5ccb77a3d0484bf85224a3c92f344fff55a989a08df7",
      x"640a73cca2aaa3175724049187b6f9fd0894d77e7e1d5b2aa91568fb79c9254a",
      x"6ede4ad60c4b093752f274e16dd0da883f498eb89d9dbd7310e2d3e14728726b",
      x"c724568cf5b4c5dc23223f602ae0bf849c853488a651ced86020ffbba38e8cc7",
      x"39197eefe6500fe2b87496e047ba101b09d2e4e450f96cd2b49c853015047934",
      x"3bb2a82cc558cf31544b85ad51e08402b9985332924b783f14542c25ccc07188",
      x"5d984a97fe4213dce3488590fc1b8971f0194c3bd903317fa032395d422abc40",
      x"4181229c8bc070f17008d0de3f2e615a4c4276eb0cfb67271eb38d0635e6ea7d",
      x"8a977e7388e1efcb644394cd80000b5a561be19273105f1324b0b35372dae0d6",
      x"a2ab27ea1f8a8c4ee6565789b6260d576cfa9aad6745f7d4c446109ab6474fcc",
      x"2abb5242ca69a9c12eabe7453e00df40977ef65b1d925b2ee821e5705a548c2d",
      x"2426fd640f51d2410bbc9c7e894f680b72d4dc729729e7e12e4fcab26a8c34e8",
      x"33362bb0b663a6a0601d11321394d9d726ad9bfc896d4dfb0d9d44e7e8619916",
      x"7e98160db520685abfd1e20b378eacb50fa0cf6315dc81f3aff7a7182be87ec4",
      x"2d9961f9897bc7f9d7646c161b96c52fd886aefe3407e9e232152bd0cb77af1e",
      x"3cd38aa12600e0adf34285d9f1066ea318be56745efd353857a1f6c4aeccd74c",
      x"6a1b262f4826d42984c07db0513343b5ea83c58bcc7f99ac90504d77d569d4f5",
      x"437caee142dea141d55950c20f0b5f0b8fb3ad12a585efd891b6c7243c9c1a71",
      x"faa0126ad1836b5fe89eb4a789852071b251ac3d18ca6c830b68e76ff6962901",
      x"b7fc6d0f336eb5a9aefe48863798aa97b1c91685bc7194ca52147a28de7db1fe",
      x"c395bc8245acf4f6844bfd73f854d5b24bccb2a70cfeeed0d9e6dcd08f29cdc9",
      x"c5a344b2ec3bb9b5daa0ad374d84e103ad4ff0d5cacd3c815cf40c4c4c6e014f",
      x"12407a5bf6c766a8028d52cc437d577bcaf808e561408827cb11b2ffdbb01f9a",
      x"dae1f8220be5f1e7a6fcfe29ba4401ead8c84a5f6d6d4d68b743958435678c53",
      x"498208fcc09e0bfc8852f0fbba0eb92afaaf4a82abb7e39ce85f87c3001a6278",
      x"6456784bd27f87a29a7c14afdcb4785d58ffb0c97430e681317b641a5ea1b587",
      x"c15fbb8b39280065d9bec722917e4243a525c926bd88e3761733744d0f32a2c5",
      x"63b3726fce4c308c21aed5a4be0b85e9b498d446332c3114cafaa956349b33fb",
      x"c0706f736850719a89485366734d7790343edb742336adc4abc164257b26ee4b",
      x"4ee119c4d697006278e0e3580d61912ebcaa03d65ad415f3b8b69762629c4580",
      x"1fb8ea0ab15aa26c4b9f59e21c891a7e1584700d3058cdd88c71139ff2f5e78c",
      x"9f2cfef2a00657675ba8edf9b4fd382ad41ce6005b478cffec8bd72aaac7dce8",
      x"bb533b750977b0d80bc1ebde81806534e1258eb169bb0c1cb936b6fa5894056d",
      x"650d4404451916f9a5f96d2d2dfe6c69ddf34eafff03effcd3006cd36203f1d3",
      x"eb74df276b5ba55191beaabb84f804226d4e398ce5abc177bf5675db0ced9656",
      x"3e75db1808e76e32651b6e9952521454c9125a928b5306ad1eb6d0b2f80ab72b",
      x"debb387a37149f7e92efc33bba00f93c0f275e3a7e01724a2d770160af803010",
      x"62c674bc47eb1e268041a7384c6a3cd7329add9de273046f9cb0ef0928d4e579",
      x"cd350e68abbd36579bb0f216585640ee87b1e2cdf9ab0518f4f5ce428e2598f5",
      x"c3db18cb3ff68aab9aa992b57094c1435771ced09c30547c78b001cc9107cee5",
      x"f291297204ee53aa4a158e8c5af6715fded4eda22c0c220270a1efd7dcf783c9",
      x"5f955bcf48cf9986a1b92bdd73b15adb75aa5181011429da4910ddf3c8b7e8c2",
      x"035e70df522cf0d6ac494641bed2e0c143cdf3e45050b0a660b1d456490e1961",
      x"a5b755271514c9d9e0d6a6bf3d39eb45e065e3ce4705f38cf362621418cc3aec",
      x"4a8019289f9907219279cab3d649b4dafdcb3dac721a99bfcecd0b946e2f5315",
      x"acf56fd0cd272d2acc87153112e80c68c7d880cfafb95a4eee2d097b9c9c1f91",
      x"45c624d86132f031601ffb967cb8fd7f4f78ebe02c3299f024b9e65f17af8a60",
      x"568dd4f83b7d27b2e63463c066daba92e47a1798efa8833d18123479ac595dc4",
      x"16fb1ba6b061ae9da02d906fc239300291f8c7d8a7179d628de666d3412fdff0",
      x"a4e07f76e7167c0fee067d6bb2aec4c365f412c8b225e7325680c1eb43dce934",
      x"c765679c7f7762f1871cfabeb47ff7dc34248828f91478deae5299de3e310539",
      x"0bb28f9546efd898b3670a2699342daa298296c403657fdd19cc7e4f7b88d0be",
      x"2ff6dfa4ff749b8939f0b1b904675f867739c7ed99f3ba7d66206383611746a6",
      x"41852fd6a981432e76af0522e22656f7e3f49424e5501a38e1fa47a6f52e2b5d",
      x"499b6cc41b974577a3bd55a6b1a12512b77a0c8cadbcfb42505e4536519577f7",
      x"87e7bebd8d22c219f5606a0369a5a97e89d5911080c70a6bd6952a50889c5ff4",
      x"6f021c37eaf50accc5a68b7057561b64bdfceabf063efa2267d7402eac21d28d",
      x"f96c64b35522941b00e9689f595b8928e1a588981b5f92225d146657e5287983",
      x"f9498f1fc13ab31a400b3bc13f753150064993c2edecc69b0560a09f8c3f5990",
      x"864b705e5b3ac64ee2745cc998685d8f2cb3f087c2efe545e5ea24fada4389c0",
      x"5f1852fc61017402daebc2ee3e0eaa71e95fcbb7de47d3eac88e3d93cf4b709d",
      x"fa8530f97926eb5f7f3e5f17b0414a89b91596dde717de391494a6da3ad48210",
      x"e261db214615c74b978afe04fa529757091e1a1a25ea96426eb7368ff63dea22",
      x"d130c496978c008c855b402955e3f4b80e9d4c4f0e5d38115681bb0c7c26a602",
      x"3337feda45ce06ac79c0722c7b3238bf61c302f6b80e7bac05a42da598cd02ca",
      x"cc5f468f9708c62de9e1ccfafe5ce7ef747fcb747c23a64db1a20ee66b827820",
      x"9cddb1f429a02b865a9e9be5f3c94653c90fbb44703908cb8672816cab437e7c",
      x"ce9387e29aef7de022a70235f0bbc54ac6375ef4a0eeb66f46b2070aff283716",
      x"86e8bea3d91700e22e6c734b9eb14e57b96922a9e166797683333549db7c73dc",
      x"4a116b58162b1cfa7a669d63dcad5e88c4884188b9b53d7ff1a243e5442fc1a1",
      x"8937eacf87cccc012f843c7cbb252a4007f669849adc437bb1fd182d24ea49a1",
      x"37aba9e891b322d410b11c94094fa5dc0734e1a9360b8b97b5fe9704efca2b7b",
      x"ea5f4a1a1c423600108f9c7211b2e63f3c83cc7dfff58100cfd1b2e96e7c52f6",
      x"2d27a2c579ba06732003c6154e05a7df52cbe602623edddb7414d06fb4c20e6c",
      x"8a80262b1a26f5da901995fb03430e18e776b88369cdb3f6012eeb15ca2331e5",
      x"d7d07e8c523e115a3a6e1085cd061d222969215dff4ddf71689bb56df5a0b8d6",
      x"dcd44609aaa7d7c7612d6ffc4ae03d476e8203d6fe07a9294c0658b6207d5e25",
      x"3bf7a4983cbc2f0db684716ed7d5259d5817b1a40982b24ff586eb77183d9a11",
      x"6fd82a1bd0aafaca0a6b7cececc7add1f42f9a9c2a856cadb49df628ceb87f31",
      x"8c5584b9bb318edf72e52c05edaa2be6d30e533414076f9c814b28384bf1ca4e",
      x"ff4a7c0131207d1f80ce0e06294fe76f8491afae57dcde9ec602ff7b534bc932",
      x"3681d490cb5476fd74466ca8ddc61805a7c319fca846d01fd06a42ce5855038c",
      x"6039a2ef9430d060ead71922aecc88f2bacc401eabcef02b53a49abcc2180d4e",
      x"758fec8aab2638b8a1e1adb3f1ba46f1f5dd63a949c891da9dcd0274f7aa089f",
      x"03cf93c4f5bf130681d0795c7567fbcbd229cc4e2f118ce8fcfe807f3fbe67cf",
      x"17f01066b9ca8499edd9759d1e44b31915e6fb884396ae7490548c7dc0d7c110",
      x"3e7ef369df575818c175a8523e295ab3e28aa91de52fb19e013c76d83e25351a",
      x"b099a9b1336718a20c39feb932964eee24546ff700db18532aebb7b3b0d85dfe",
      x"8677834f9c54c532fe052b9cabc002aa2d84be4bc0063a98fe47a21d3211cc45",
      x"d11122ce632abeb52354f5ce22c18aad8775146ac56125bd6fc1a2850626a91b",
      x"60819def0e78bd2d5038d3208e804d36bacd5059fa0ffccc40d288697063fc4b",
      x"44766f82d671c1bcd93faa89831aa51440ceeeaa3528b500a727f6ed354a2e58",
      x"faf4eb367ed9f27f6cdb1bad0630d3c6d3097071c51d55d504059be8ef979e62",
      x"cc28043cd07441632c97b4e02dca80fd4d50d8915a810d85865264905c50c934",
      x"fae1527b9eec142caf41ff92ba27702a574d665e1c025d8316086c6c69a507ca",
      x"020676a045d37205b58f62e24598c0c109c9aee6c03355a24a1e20bcec019d7a",
      x"0c35fd60d336f880adee00687da519aede00f2b676c3dbf47ad8d0fdec0816ec",
      x"8896e457e6d2758381365f3cccb6e661d19610a482bf81b6474db8557cf600c7",
      x"1595e6deb2828a9e96883932e1ea0f071b78f25ac6a62ab2e5a25629c2b9e3f0",
      x"abf730706927d814a232523dee110f62d9f0722c2decdb945503f6e62e386f66",
      x"4d83b40106a09b9ce74529d735bedfa995011c1b588d330b3bb56dee34fc89bd",
      x"f955ad50dde84813d46e961c71b6abdcb797e56707de124c94bfb096ddcabe9f",
      x"40859024e595a6f8e7b9e5baf23fd493a46f4ae6cd6774497446834d3b4f6b76",
      x"6c71b5b4311362e68a753f08a6c042f523a0e993d939b864b5eadcfcaf16100d",
      x"1260e7cec31a3f328e1936fbeb45e0fe5345973587d6bed507fab05ae5163891",
      x"d4f37aa5666733d106c0e4b0fb050d67ce7aa6c7bf0f62107ff955810a32f7cc",
      x"14316b35bd5876210c26772519287dc1abb0ef24aeaeaa7f5d4823f2d589706b",
      x"b35f9c57c4a3ce255e25bdcb2ad0bcf4a3484a5d5646f4dcc7d1f1e0b07556f1",
      x"75f38a8440945af746212f2ddac26742a46327aa73775493a77f51a008e1c04e",
      x"def0be6f5ef88cc6779d53833a467e83249cf99c10b346be72b2cd6c0b8f734d",
      x"79ae4bd0118afa441534ade6e9c35d6f7f81e09c56fba80e46969b508e5755cb",
      x"8f201972d8e1c7533dd196296b6fedf969cff2ac5b00ed000b0f7be6fe5d9578",
      x"fe6b52abbba1f1874674cf6d00c4c928ae5aff613540bc892a5112528a694aef",
      x"46c627edde4e1855bf9790e181eed23bdfae01d4c9f5e0725223201cf7fb2f71",
      x"d8ab6ff19eb590383d6512ff05040f8ff0283cfe546c32c2b414641722ca1141",
      x"658dfa503302e7a07a76946917f60d52b0ce08810a1b2304c107bd36a8668fef",
      x"51e5b11dead742e39c1501d057862b50c8d98133a6add75f5580e949bcd249f3",
      x"e057911ef1e09fb5fc371815bb51c62d2b544dc8e80961426fdf6190bec4831c",
      x"e0b760f96cbbdbb2466b5db89f8bb7804d6d5b657dec00961fca5881654a443e",
      x"bc418505c011f9ed7e9b5348f9933ca9002c8a6f39599ffbc620034d9811da4c",
      x"7b9b5b721f8f288f560ecf53075b316b0e32f25b1e7dc8d022ba7e1e4e4f4ff7",
      x"aa81dd9afded33cdd683e9c5fdc81f3eed0002f85f7c7f343c6c1e13afe3569d",
      x"bb7b3d49a6d0bc72299fd922d1cf31d97ca61fd49a2d51a9db8be265163bff0a",
      x"84b55f62e45128a4931cc2a35d2e34f2e8e89a61940eb7c14600fee0cf053081",
      x"54af75e17985076b2ae0b7fc7eb6ead4944239be9ecdaa7866fb229e3b8e88a2",
      x"ca8cc2cef51a771653379c46bb63283120b95c97f453876e71a5cb5927f9af5b",
      x"29d74bb6b4fccd6cd303fa4656566d2c70402f2f2a02eb6935107dd9a99392c6",
      x"d0de7e38cf99944e7b2a8ee99af5d2f0d5d84488abaa13f87f505782af9e6c24",
      x"f86db2a1f31e67f2a155591b1010498be16a674dbffd46b9240fb17181add12c",
      x"0fdcb8a0247b99f01830d3b5fcbb4ec97a88a8fb5a83f8f33ad43e1684f85d63",
      x"fa5c9c646f15a8797a9fd877fb9b1911b6aa8e313b6bb50af987527043ec0706",
      x"382d6fa65dc92677089f1590fa9e610c8db095e8402d98132c6badc1fcc6404e",
      x"715b851709a66c0292968964ef1ae5f9102ecc462753a0a3a915c653742efa4c",
      x"5422ce2e0128b67956239e219a38993f882a436b79b94e63929faec1f0afd021",
      x"b918df7d41c51c541762168a00923218d7fc5f0583cf4fc8130cdf557f9621b2",
      x"e429c69ec985535cb2d8688f434af119f2c828183c128e38be9ff641ff0b06f2",
      x"916cafc074e3858536f23c6d1c1d6693b3631eb91aa196d1da76641666940b94",
      x"2b500358958502caacf00e1de97c5728b748371080a8170b217d2bbf6cff5ea7",
      x"53b2a3e636f89f1f800b9528fcd5aa2f97d57e838b6e9812c524acf39d4caed2",
      x"1c9efa849e8f065cd02479a288e3b36f5dd26d7f711aa08e4c198fd4f0c75472",
      x"c52277e4a36109e382e4a9ca9131f33db62cbcafae4ee5bcf143e62bcefd18c0",
      x"7997f26bd293675c91b95cbd16f249ace313d536ec7f683d141352c85e62511d",
      x"67cdd4133cf021207076ec337fb0e2b359933b07f493e37e3f6e49c6d94670db",
      x"94f94eaedc69d0bed11f2052074c0c930d29baa0f3f6147d44e042238b0fa499",
      x"bf0508519d744f1779a6b740ac9ec86e6b830f558216a96e9e3b634f749f74d0",
      x"12cbc114bc2e644b933c3d7de0b28f95b030981d5f5be6d0ad812c7659b53ea4",
      x"1c8b6140504e25ef99af49779a0554485dd6340433194c75860200b5635fb5ed",
      x"3b25f53ad1df2b288e59c869339ba9cad6369b7f4496f6817ff2f1782769704b",
      x"a9bfcfd877d39423a8b540ace31bce489a7a50be21c3be8d12dbbe13e68121d2",
      x"13892f603eb17958157fbfcae90b2cce44ce753fc6f963d96c90c1442d4c230b",
      x"5e35fd6d0430fce5d67f03ccad9264f0d6774ddb7d975e14dce68aa486bb7bc6",
      x"33c53e97a71314128cc642dcfa0605024a45a209004d749c5cb41ab4eff8648c",
      x"89b2d9fcc35013f33ec28d2e6a787c0c12f589973d94c35a5fb03ccfc2f23238",
      x"79a77f9b5dfbc1ea43008ddae6c3c9ad3c1aaf88f7978db9372dc243326b69cf",
      x"3aaceb45f7ffb40ded04938c422aaca930ae8b0aa94f14f8baa545471f43f3e1",
      x"903c26173417b6cd631673ac949b02cbbf04e99e31912bb59654cedf52d1c963",
      x"7fc42431bc141f635135fcaec683c517f9f18a8e9ad2be68a44f16e8da40d178",
      x"d59cbd50b3576e4ed94859921d13cc7da86630ea78bdde64f64d9bea015959d4",
      x"a39108b457aa2632e8c234bb19fc26d3b43ccf9b5660836c1501f9ae9540db0e",
      x"d0a41e59387839fe4fe1c57bcd11e1e28be6948a36e99e6d71bcc3ac3749be09",
      x"7f2774ec1a03885a8ab4976e3916d0d169cc67f61288a86e072dad77acffaa12",
      x"8233688a336818e9ad6cd666b840eb23cec691d207d4448a045c7d3624050f6e",
      x"bc6a9b5bed9790aa3c14c1cfb1d6ac052d9dc046c671975ca4feeee733bb5aa7",
      x"84e2e8df8c778fc37c0cfeb1a6eb5e0315e41afc3ac780e639e355d2f36cbeeb",
      x"d7b1f0c54f8d71edb65c060abee3af35ed621a477dd226ba67aeccb42fcc8a6a",
      x"c3a3efd0d74d989269ffc2f39555fd3e13a1aea6ffcbf7de6908ac5c2e8fd529",
      x"726fe653fbd06ec68bf8f5b9a3c070f0fca61ac5efefb7705d06b7d6a06c023f",
      x"b61d10881d4f846549d9a720e37bc95e9d4d817a616f34b180ed146698a92b05",
      x"f3602db73cbd764f1ac3002a85329673373fa90ad5d63698432c1d62a0668204",
      x"0aeeb9aecf815f15e49f1f4bb1692904414cc1d6f18c9410dab92ce0352ced56",
      x"f5ddedc3d489210b784e452cba8ff49781b52dc3fa79632b030446e3b64e5dab",
      x"0ec76a6534ad9c433a13e144de12d1036fa51b9c72bf02e27f0a5b8e43542b06",
      x"92b5b5a519879310cdb6fb3228ad65395475a9a9a3ad1670a07987b72a643da5",
      x"1717b6d4cf900003cd94653d4c1e7d7be27ec7432e3c7acd8c0f444c170d0b1c",
      x"6d0372580700959e90be4d7904a0f39bc81f900e665e51cc17e27c44336afe56",
      x"d5609abb817dc7616b7cda8d5d8c3c4f35411dbe0d75af8ba25f377ca1e550b4",
      x"06a98531866824815a6ed8b457603a4a75cb7f79ea11a96ae3b9ac5c36e7138f",
      x"6081143b4db30a1f3037a8c0ba3fbbcd9ea7cf60907c7bd49ac0a1430e8eb774",
      x"d1bfd4f6b2655fe67801383a06b2b4aa185a8bcbbd15cf6153967da1511d03a4",
      x"e583a59241bf994834da8835116b2c76c754acd050fcb83ec1c840c1c603c8c2",
      x"9f07d1a7b59db582fddbb4b7487491e53c71c6c6eb43bbbf83678a091473cc05",
      x"feb88b23c6070f789b8198e7a5973d93ac62ca237588cbd4bfb332764006bde5",
      x"11ec68dd9edf343ed594d1cfd5ae66d88dd5db0de56e73c8efa57abe70df27c9",
      x"d813c1cd9b3ea5b87524162ac7eb7ed16286002a7f2c6da29ac4f774fa53bdd7"
    ),
    (
      x"581a7e407d6e6548cc1d70f3e590a3e4e9e5c850ebd69bc33d455a93db1ccb1e",
      x"2d6d0101426a455ecb67a8040e5e1c9f0668b7b5df4867bebb05eb1aa2c1d923",
      x"e6b1c639d17ad5daed89a68618faacd2085eb3cce3097f94de9de4d7d3a5cfef",
      x"123511d5b15cde3d51a53913c717b69eac1774d09814c636bc777ed3fe64d387",
      x"74a2a904707103c2d6b17bf2930eef2139068540c2994e78d62b2ab37f317d83",
      x"ded3576bffd84958f752ead2df1da8cade977c16ca9acf3daa5ba867cd1a3a49",
      x"bad95a8e6ade316ef02c5bffed8703111003505a579558ea0fc622fb2d2e3748",
      x"c799ada835f65cdc51d4eacdc6893259a244f20bf0bb13997e963b8cfa0ce729",
      x"6b1caee826cc843988692bc0b921063bf91107b0e1b8740f8312f1c8a27ec94f",
      x"4cd115f06b59335a41f11d7dc99514628ff40df74dee2fb95f007022266786fe",
      x"fd0385c8cfc50bcbcdaec197e6cfe05debfb0af601259f0e68887163bc20a288",
      x"258e0e2cbacd6df76704102f0215315901b04d4ccbe7dd9d0c57b1aa8aefefba",
      x"5d8425ad8c903c164f9f52bb9544d31bd3949f7ca990093b7ffe043d3b954a6f",
      x"b2e291242ce1a9457b0e0ab0fbd18c68e97bfb892c85e41e467d304741ecae57",
      x"c7f94b47f3b4a4e0fcd134e4d6624490a4a0243e219c02bbebfc094e573bde62",
      x"7dfc516d8ad069a543cb1d8ccbe19d9731ee128f0f4dd262f3e9b5fdf3fe9f0e",
      x"4bd2acbb0a0703bf824bf68c4851255a0a0abada10bd8aca3a785f3f5cd34f22",
      x"6337d4211a2323b987d8687b66b0bb5c00c98ef2bc61ed33457e3c75c5a5435b",
      x"73bdb7b658ff2330fffa79783017f81403988b37a6b2745b8a6cce38dd065f45",
      x"7b71f91e2e5b6b840f12b149b099c0be2cf13bcd31af3dfcc053742803b7a2c3",
      x"2737133d23687f7be10d47bb5152148b2d77cc03a161f89fc4cf71a16a752504",
      x"0024c157ccd4c9bec888f3278628a86c6fd84c59893b11bc906d1f10bde4b85d",
      x"2f60617c282e2f7978f12cdc23aa6c412b13739e7090daca15cb2072151f0048",
      x"b96f50daafde050edb17c7e9947337783e13875791cc67bbb671c58d060e2d83",
      x"4762f2fd740f8d572f29f94ab003bc43c6776ff79b17b17cf69b3785c55f34a7",
      x"c96297aa4ff900d8616aa99a81e7d636840cca5f800f51b52d28b01dd3440c84",
      x"0802a6bbdb19af7dd406e7e5284c7058bda13268c4a2b14e004c6905c255505c",
      x"57ddb795da0a40c53162915b54f8087cf2658c6e1af74cf318e6669692f25243",
      x"0a563d3fef1d0d7e1fc2fc42c9c1fcb240c7fd66c6b616eac767442880a078a1",
      x"8114f96db31ff387df89029c8dee8ff35ed6174bf3e749979dde628e1c1fd0f7",
      x"7623bc47e9b23566c2494584a0b5d7f4e87f52c7d23023191da0867b03629bb7",
      x"41b08117eb1d57c76a876a27f3f58e64741b986a32f32ec1f8e9d60859f70b77",
      x"e8fd8c3d33c506196664c7801766cc1b6b80b02c435bd59fe2078887741ccf81",
      x"c42d7cbe1be676efba9d1f2f838fad11a9a6b6f0a832c4f2e5a31f6bc5ff616b",
      x"31f8498b4d8fc196a63e01279c73e4224776ade77020a743efa45e39e7063aa9",
      x"5535e2be194bc2bffcd1b690e0a18a6c0d935d299052ae4648696bce2dc0bd9d",
      x"0fa2ce383bd6649c6da0019a05e95f42e344b00c5b62d74ef94d2bf9573c0ad9",
      x"da1e127c95f847236bdeca5c0709ff96f50455903b0327541a3642cbe7c9c3f0",
      x"147f9d5bacfd3bcd5f598d81392809978d1d92645500a02177b76d31161b5579",
      x"871ba00c26b0956af898a0588a1b275c441f8b530333818fa7f5e71e41e80593",
      x"3b26f576ed531a0f655a4f3abe4ef053dca5a9c7d1f678d897f189ba73863525",
      x"10810d026a586a20737964157b285384f7c2d408a52b1a0b15a066ad37bd7de6",
      x"0b7e138ab2df7d942f8df558655a24ec03ce3e579013f90a34c02580e2f9828e",
      x"8a4dcdc475a046e76f0caa006986bcfaa8fa466669eca987c35c7275a8145e3d",
      x"121876e5708b0c6d2eae9b949a9d6dc87ab740908312faefdec6ac5c80a65c65",
      x"33aaf5292faf1395d853e2bc5b4abcb557116bd7708d0d1d97c2b4d9c4f7c3b2",
      x"63e094fe7e9194fb7674453fc2d42e32cf199da496cbcc55ed127958b15d2ea7",
      x"dac1c6cf0af2543f12bf23ba172f6564fa7d4fe804eeda3f82536f5e00aeecac",
      x"270af88943bb12b6eb50f7a44b12897325e8d41b423ffb1bcc5aae004e7b61c9",
      x"d162b01aae6ba4d240290a2db22f09d7e545fba06641d0517ffa71e6cda34484",
      x"1a82fbab5bc1772f755cbcd782514c21f59960e73375b20a91ef0d31330455ed",
      x"2de35a09285ba4682e2a964f0288fe217da5566d4488c25f6a85047583f106d0",
      x"082f56e36a6f68e28a98c3a1af65b70985e69d8a65e07df2867edcc561b393e2",
      x"a0f2031ef811719f7cd7272dea678b44a11921c4ccf54b565ddba664b8d17403",
      x"14730598a507095a56cde297382f6c37c12c6081ec415e638b7eba6c9f7f50a2",
      x"7e85007d5aa68c5645726255de7b88475c6d1bc84a98dc1fc8fa880513d8dba1",
      x"288cc6824b2d1711d5189ba47ca614ed119bdb8d0e0cd9d38d6d08462d992477",
      x"ad6e8efb53be72e6d815e76a45e665fd57f585f543876fc814ac80455a4bdf9f",
      x"249b1f86481a28fb28960a4e453be2028227a8c192ceba97b40da5eb91970af9",
      x"c18f1f246fba03984e39a1c3fa69371a2f6dd8d443187cbff701773b3163646f",
      x"40dc66c55c38929d6b36b22477ec2918a39c9ed64b11747e91fd90721901c045",
      x"86e7b71e5c6f46c523ab81842217cad06ee12a99cd604e40969fb83d3644231a",
      x"2a1198de9c7e252c326fb203c2bc260a6298df965e5ab6a52e5a1095f99fc216",
      x"b62da41decbe7663e2d8144c1e4f7f7438bfee31ad7992ea6221c6c526ed74ca",
      x"dc3a7b327ea662912a2e0d328b47176f5ebd891471206af581c98c618811bf23",
      x"2391679f38d3b53470f55520922c3d93841dce393ce4fa539b2e81e10e678846",
      x"b9ddb4289db701e9776d476bb6b0a1e6245f9aee4e36ad097c6f6d9cd57045d9",
      x"99d81d5881f3b7bddb846f6a87a36956cf5fab99dba2d5108befc933b90036dc",
      x"5dea902c3469bbf626d1259265bca97bfeb940ccb3eebfb0d26ad7f4c6bb1f78",
      x"a68669aad7fd2210298d7f11e01f58f60f9be521b9be7bbbadaafdb1a1134e01",
      x"179554f365bba5b962ea7676fee522359151bb7d9fd5cdc86226fe7b4abc0d14",
      x"f2636270aed98709c850e5fdc9cc60ea40fe7841b33af91a35c95c18a4a512fd",
      x"e3077a45bd89da317e1573c86af6e9b6de465864a8fe96819e2bff56c430c45e",
      x"469cd54fc570c074f3b700c555dda121abd76fe9ef2e6badd41f8f6ba316b122",
      x"06f6f8c72a2665765818080154ac0531e8e92a5bcdc0fb8fdf17c5246f88ffc4",
      x"d57e0e20a79a527a8cb8da3a1b9a40fe5a2a6f5a80238e617f7cf6201b94a4ce",
      x"70f3d8e70546e2e8c7ad56920ad798fd9cf1f53970b4cfa2e1dc5703f85c5347",
      x"bcf656da6f623e7c9e74dcc295077f70bcd2765003fbdb51b17fc8b2e4c24816",
      x"e8806463b3965d27fcc3a7008c44b8d764d72bd796d775fe0c7115a1480de6c9",
      x"497958b94d0c0f17c787264e1e06fa82241ab5ab8c8c69c08999dba89e58d480",
      x"8dd321d6e9f12ff2cd9e75b153c7fe3b2ee75223f9d139f9afd799f2195385c9",
      x"985bc9f93b3503837a52dbcc227ccfc2266cffbfee478bf6510843955d5beed8",
      x"92da7984fb8c18c930883aecdabc31d25eb057b11b9c58590803809b1e3aede7",
      x"064bb0e5fe692f809880965234e60b1f01eb695b04447babb1fa721c640dcfd1",
      x"4aa0ebfefae873204a8b20e0701f660c715615c42bec6af3b7b1ce3aa6a56080",
      x"7c849124aa9bacb93b5a5a30d5f91f893c8086ad1527ac21a1579ed7bc9bf34a",
      x"ec8fc9e628e2cd76e4a7988e0ca9307a26f02236a7e91e9da9257db310fbe96c",
      x"8acf39bf2923efb270d74a7e2406aee86f593e5cb0240b749b801db1d8d5ec39",
      x"6808789ce20bc6ad762c1783c3496b76559b82d7e20de556ed174f4ba5e77788",
      x"10167aac350cc75c2f252d378bada1c2abdf6940dbfba52dea6e9314e0b9a3c9",
      x"d92266e1692287fae50829b01f4aada935e5e2b5211de15e459508b1d4994b11",
      x"97648e670f6fcc2d3113ad46e66831112d884870d5053384dd37e167cb23b904",
      x"aba8fb939faf783b7cb16173d1a2b9189a157d337b429f32c693271b38f6b8d4",
      x"16e7629764bc17baa3609ac47c180e7b0918ea353aff9f86c47c686922097177",
      x"482be2efcd64e734881949b691e98f027ee39d73a0ebbb637affb9aa735a8953",
      x"7508e05198ece510c67ce14485460f9b63e518ec9d84cc806f160023e34fdeaf",
      x"e0a151f501c4700c20f6b91a44e281c789f2ea4ff2d90327560ce0e51856ae92",
      x"20a27321b76c23f7f81f471f899b691bbe1ef285d385d157d0e7e655202ea9ee",
      x"0cc30db4c402012bbc030b629d141418ce84d3465fcf3e8a9135eb7229ff730d",
      x"b042be76e305dc1bf8650f5f04e1554e381d297356ddfedbd26f6516fbc9a493",
      x"d810ead8319fcaa4016f11b640efa14f792883ad7e65a5bf2a333e89cd3a0902",
      x"2d9fa9f9721502949e904a0c37a6aec3f07257101b7ac8e77f290a12bc01c8bc",
      x"186ce51b998ff827974d3ecb88cc922bae9d949229634375ba3384d52cc36e6f",
      x"6fd418a949b93c675f6c02a8d86bd79ef4439ff42f1befd48f3242242ac23636",
      x"11d2a2b0b0be693b551fce98a03d86af3c0c105f753d16571046d2980e0a2e8c",
      x"9c5a12f1b904de502e2b9d80162e9498db4299c1944e038b1e811e1178f9aab4",
      x"305b047eb846dab9489d7e9b3f2ff2e18ad010cba9d8d582eab5cf0d294026fa",
      x"8e4e6c50b48401441745a54c685c29f6a4bca92e78ff7640c3a2acdfe6cdeda7",
      x"e2f572ef8cba04a1d3d3f1e64f2e11e9cbaea876a331bb734cee28f708d1d300",
      x"c24bdbd19db1aac4356a6d079200462327e260d84db6791674826b2f137a8d30",
      x"370563115b7f1f48758582056ada1e7d2c76a7c1eb1fe024cb9d262471eb58c0",
      x"871b9a45268fa6edc07dc8ddeda56c4e13dd27178c7a645d549bc48d547ffb0c",
      x"e68082144ae65c9b2bf0899344bc9a364b0e25e5532f93de425386346cafa632",
      x"3435f8f083093920a4d80ade73d8bb9e1afe30d19ca3dc8cd52fa4555440b6fd",
      x"689b7ceb5c39549e036217f6f1ad3080b0f907e3a17b4ad110cfe6bd2f2da30b",
      x"8f0b91af059490ddb1b93ed2373ec3162cd8a320e3cb88159888aab87e564cb9",
      x"524a8faaac0ad116af7ccc9f6f396ca5f9544155eca013eafefd2b98bf1e7eb6",
      x"053c06e5acb64b8d171b804fda5eaaf1d35ddc54d9895039912331d0f6c47c1e",
      x"abc38f96ce9305640dbe4f76dfd273e6941a8efb8e1dcf9ca7f18b9aad3a8586",
      x"a5a9132bfca9cde2ca640429a0e5efdd9b75de7cb79b294483a414fb0c35df3b",
      x"82e22099bd65aaf8135f45f06750b39ec31cf7756ac0ad7be42bb3773c13bef1",
      x"a174561dcf4563039e8018b3465feae4f4dcebe79e197ff4a1f5cebcd8206e94",
      x"7d2828ca50b1bb78f8b57b666b19f388414132f390b3f31030cb9b6ab2f917b3",
      x"ca44ed3b5d4469d388b4ef0f24a5054af03173943e3fddd6aacaa9831f9c1a16",
      x"f3343a8a118d9719e8cd2177ada193aedcc0e2b44b89862898cbd4b42c7b3a02",
      x"daa84be59cf3a681351687dc70c8ae60e66c289b5c8c9bc39698241985de5452",
      x"d15c4ca0b0280ab209e6f06b646d75d74cd03b1207aa11bbdacae3b96fa04c2a",
      x"55c3d5a4d45194d3342fe372c220ac55a5ffb9bdaebbf7e00496d2ab39eaa082",
      x"e96528632e3dea25059677afece4fc074ebeb0d2aec16873704e2191347ce7bd",
      x"c7a0508bd4c04aadd1d176a1e2459e8057e9bcee059f0221f5aa395133495e63",
      x"1fcc5ccd6c297f23865f7879501e6e3852849ef54113bd8a841f2606e3b559e4",
      x"71380fb2bcb222ceb8c8774460d4c0bc845365bb028bfbbf85ed838def631087",
      x"cb2f33f4357773a4c8dd0cb5be260b60c67b56da17a347fdd62af8b631ace89d",
      x"9592bb27c25c01a6c27afbcc41829bf429c0c8c11f58a55b82affeac4efc9382",
      x"98e5f51fdf49d021370bf9d1a75290ae1ce90e0a29e59c75bbc81460338cacc9",
      x"3be043055ee9a786673e7b54685bb535ecae1ad52d2301b6730645467ba95f0b",
      x"0bff89f8554cdc29035e204dab4816f2ea1e0b1b1ae4a4de7233899a675b7221",
      x"1001dc8692f59c875883fd635dd069aad8769bb69833441c2ee0126eb6900b9b",
      x"7a3b7ccf910660343f05f27fb16930bb504783a9cdbf635bb308a839c04fe5b0",
      x"486faa6e8dfadbb35dbf89de772c720bfeb4a334608d7f1d3f4dfcb96917070e",
      x"c83ec48e27251039cf4da5e75b69caeb915ca230ab39a2d6b7a1068c0bc360f7",
      x"8eedf8e478742a56f7b67ab5b29cd4b8943a697901c379a8da567e0f643514bd",
      x"e499ea84b1ab965e7790738af10a135d0b7d86568d56174773eba5afc7a24858",
      x"a512740de32f292a7a320897ec78e49df62976705668902194258f0cf17600d2",
      x"f7135f827f44368e25e52642c42d97f4746734b4db41dec084f31b1e22e4928c",
      x"622de5f5507e5a1b56ca3b7e844b7578ccf3d3cd6147a6e6a0d8c3c9a63ec750",
      x"5c0005093db6ad361f283e5b962bd1a8548aa45e9144c9e7e01f92916810b473",
      x"3c046cac503963400f34442206d24d8f77f3d72ca64bdebd8b040dd13a034b93",
      x"13d12f35fd9f4209b9e7248cca5839df96a55ca0550364fcb34c15b09a7cb291",
      x"43f596601a71528cba848aff5fa66fbf8c7199c5fc5e8d9be24db358b55626f4",
      x"73d1eae55d86b8357264136eba00f29bf75af7e961584f42f26aed0ebdaee907",
      x"a943773cd3f5f6f51a6ceedafd07f73a50d13a23847d4d17dd9ae06790bccf53",
      x"00130147fef7afbb658916eb5f14e48df39026c191f0a25f1b86646849f5af5c",
      x"8baeb7b9cc127b868d55d12bcb95c7a6b4dd3d5b4e3f762d41b0b5571c900a8a",
      x"c026d9b256f24f1e47d73aaaaabb695e625a3b0279b2b7f57ee6441c3ad4d315",
      x"eb07530e94ec07081312ed196caf1243db5e7ae4dc3c3e7b3867bba99b14f3b5",
      x"d643807639125ecd93b25c72565b253c060cc2e06a1ac1a70cac5b79f1f17966",
      x"b5d05959e9cfab9ad52d88846a5846d480b559eb85c95ea8bc52c6cae8d00125",
      x"941eb99454e17efe071022772cb62ea086604b6c4c9334561e117ecedfbb7976",
      x"5644092d9a46f7f692502a3d54459c72ed2618e85b5fa447c00ffe5682b6da04",
      x"bfde1bf7dcef0336faa63c4972dc4c2ec5819d528c4017ced83a583dee7329ea",
      x"308d5bb31c2de8b244a7b20d2090fe0ee6787adbec702edadda8815be64dbff7",
      x"aaa2618f33d63cb52a4e33357d6811bbeb77c9fa8bc142a363ff0995f97a7dfb",
      x"fe8134296e1605c1e952b257b3e20966557b413bbec6ba281550d8b6f5e7c2e2",
      x"7207b930c04725470c66056de9516aa91a4b10cf038216b06e62686bcbe3865a",
      x"bcdd04a9efe0ef943e4e65b4a73ea32d0cc9a76c7e1d33f88e436400d3810815",
      x"b9baef7b397b1d57bdda2a8b035e10ada4fb109ec87ab0215651728939521d77",
      x"cd6aaa9fd8932c63e2fc9ebbf32b119853aba16c87de970d5b38df1a2056b454",
      x"3f9d257094a68a4adf0e2c4bc69c129bfa70adc411100cf48094789d311d8494",
      x"8298a1cfa5ad41cccdbedfe41342253b934fb09fd4009f266233479cb310935d",
      x"f809f3fec4e6d2073beb3d36fa6b93ad1248a4aa6c2951f7f7e0a297e50652bc",
      x"efb1f8660958328e0d731f552f620702d23d0fe27dcbd583aff831e64f486c5a",
      x"ccf34282055dcb782bf066732f018edc9615e9f0648489b1a1e137ee3c0ae536",
      x"3b331719a072d97832683c6f0aa2ff0e38f256e4557b7738200a27f46d3a0ca2",
      x"2da14cd84a8d73206b0dd9f4bb9857a0fbabdf5b1773bf714aa3569cdcc78a48",
      x"ead520d3f5e47fc2e3ba7e47ecd27444175c8d6f35d4380b941b6ee2f54ea06a",
      x"89a637cbccb4ffa40504cd8dca647e468e35d30dbc654b4f88ed19e364d3d017",
      x"3a66c1008f5055b38326cb63b73f6f03da9db6ac4a00f6caad27d79e5eea0744",
      x"ab9682245e3105df2c22f6e5962e179152c33132622f2ab48dfa3161d4bd72da",
      x"7b7d5fa3b731ece4dc2835074c0024b7af7e3970bad021b57fdd1420f2abf100",
      x"ed1348bc48e219b1894e324dfa48998f1185404e99cd20f416cf1d7da19e96d9",
      x"47af49549b08c6e7132bb6a3525c232b36f52461e0dd5a6771e8de664cf788d1",
      x"256f4612245ef2e043f4465d77b7ef42bdae1bceb6a7a48427c38095230d0301",
      x"9744f6f4084d0c462c0c5a5a350f26e0c02ed65df094108adc8cc7eb0dab08e3",
      x"499187b2ee2062e9a9e9ebbdab9cb007837209aa3d4132ca55ff4cdbf8a40024",
      x"b571f7e906378ff62d93ca77515d5254c35b9f0de5cd84fa28bfefc377d6b3b6",
      x"a99a5fbd745bb16574203868029293b40ec7dd25597b4b1069d85944b63aeb09",
      x"db1ecef73bfb43ac870bddd27122be7cf539c527cf4b5eb1c4d919598b23f9a5",
      x"41a630370441493cd32b18dc73e8afb0f220066dceab464c5853951e2558b8a2",
      x"c53bbe658f0d4e681ec7b2cce4a005577a2bc1ab13488033431b41c419187f56",
      x"5ab2724841425c2e28dc05d77ab43366f8316ce1f656d8914018664c01376e2a",
      x"92dd2769c83bf90059700a43ac6af053e715ea10655e53a321c5ee9c81a2e402",
      x"715c47d6922687f048dc0d7e8738ef29d8c143151481b5b648b45117246d62ca",
      x"fa76ff2fa59fc6ebad9e41cfe3fffccbb7eb2d82adf326badcae71030299becc",
      x"eb04cabc686665311be91fa68724f2bf80e90a396c88056f5e20b308c4adc270",
      x"ac356b1de82df86124986202386690457d6fe7ff1a8b1a1c172c01a8dccb42f8",
      x"52b57cb6c0408d58a45537383b9aeed71b14c26cc8890e46b6a4b3c9e3fb7614",
      x"bcbee83f9560a5724a552e5b9b22d9472766611dafd57002b317bd402c2288d2",
      x"cdc53d4b3577a29b4b4f2e5a42acb295b095e53fcebc5d5f1ecf26f34eefbacf",
      x"5d6ac02d311beb7561147ecb5d6388e20da4d6bc2e4caae4db7e5204a15a863f",
      x"f85052fe863fa1a98f1e1204e9a5c7d24ee96a3f5d9ad4ea6e670cdb97fe2a78",
      x"cd31e500ea69fc22be8cd2eb86c55709168b6e4a4b3c393341d4ec5369c653d4",
      x"a0c2b4645db3014af840430f59b6f0da8619efa3808d9fca17486a5c1c5be949",
      x"a2b307da7051105ca5d6c2f8b9d90061f8267379aaee38696c7dc84f3e829596",
      x"58f2fc3c9069dccd91808e6cf8ab4bcf63a3039a2278208cddc4c33a0b9bab5b",
      x"8c6b4192673038d4a738378b33e5f893cf4a5713e6c670815bd52e6ff10033d9",
      x"59a70889e4f6ba85ef790203f083ca79fd172a8f2c4d57f0c22c8561def215f5",
      x"4716fbef8b622a39d0c487afb6947f60de126f2c43a4b54e2440cb6bae6e544b",
      x"c3a550448e6d4f0ec35b4fae4887ee994e94e745de12aa0c3cafa2ea6c443656",
      x"605408692c649d0d4092fe53c59b8615224ab435969a30e8b8348642ea1706e2",
      x"8a72f525afbc6e609281128b45e70ebd244935bf6176491275c092636df858dc",
      x"01da4f459363deee36971653e3c19d2684901b486fe9734ae55a01257754e2c2",
      x"ee2ae3c5f085fd3f727287dcc046f9759b3c17e8ad05c8f8f1e7e03ac0984b0e",
      x"f80637c98574c1dc798c5218a8ad4eac8deefcedd8aa639f8fc627a12910961c",
      x"eb82d3ea04e329e362079872a8a7b7f11e3a79699182e04cee4b7f0a80f925c6",
      x"3bd671bbd3473dc07c092e54c9136a20ad394f87900b2b9496d6807b9be2d93a",
      x"2ee496f56d6536ed96013d49ac83cd12448afd1414ebbaa5237dfec95c3950c4",
      x"78af237dff856d35c66e0074b7a71e999ea9c5e12ec19d5aef9c4e8ada7b6893",
      x"72340cc5791ec9c17a05637103417d9e754835e0e77335d5e6e80f9b0f310b5a",
      x"60d33a140692c501f85e177439e4c0766bfe13fd7efd2897c3ded91c50306fd7",
      x"f3dbf54d9646fb7c3efc50780b7bba748f71a542a33b92fabb8a9b23926e99a3",
      x"b18f5054d362cdbfa8aa6fe68a6c9ce0a80848b868c3c36eaf3bd47f27da0162",
      x"4b919c26356f8f4122ec4b87de722111c76d32ee06562278b9f3c0fd7677b68b",
      x"0cbdb1ee6e8a94cd44045a07f9553e97764f1b3e3d4ed1cd294cbea4164ec353",
      x"108cfa028787504018b20b96fef7bc4340593df4b5e26d37af9a610c8a99473d",
      x"0ee116e35386a65d422ac3255375af71acc26e3dc1c8b666ac46931ee5d3182e",
      x"e468b6868175fe00d99b15f1f7bdb7079af04b78478028dc82220fd8abbda03b",
      x"47ac63829794f9de9102f1fd8d69abe35b54203afedd7c5ebd5d7584be542107",
      x"13d88733dcbaf9827e0ef11e4dc8ac039e0ee3ffb551a3bdfb20817669847150",
      x"0adafef14726579258b16779deee353188c2ff9159fd986ba7db84a2f40ff2c5",
      x"7c842538876dc5efdcd4fcfd434331fdeccf13c5cecce63eb76c6c858b6a5388",
      x"1741ca916fb6c65f27a16032a8065a7263fb4377b101c5f30ec8052912a8b690",
      x"6e3e97599a2d031f0c65673e6b14a5067e44f8bfa5d71ace5097c4060488bc1d",
      x"1da9c41cebfd2731adcb889f6d751bb80c9b40a078b6dad8261163eddf4ef426",
      x"74f0236d0f5d8cc196d982dfe643e741163eb45d76aebaac634a6b71ec69f9e2",
      x"fa713ef0202ee4da9b18a9cd85321f0db52d43c6671acd4c82de8e183923bba3",
      x"7cdbce6a80a4ed5a10f7848b3dd524bd727e646e40b93e10d2f8edde93a287d0",
      x"57817c0bb665a02e07d5cec1df759bbfbe0363b4312245447b6cdee78d0d71d5",
      x"a63d63bbaf095270ef399a07501fa1f8baf514e62fb3f214c347c1a4d7b9cb9d",
      x"7b5c3d8e16509596d3c400fd0b75672d43888e5200d750297da5d011f64ad7ac",
      x"608d18cb31803e46b6e2c15dd1fd4c465093d732acc61df8a4195c5c9875e1f0",
      x"a30c7639d2c6a744a35013747a61a204b0dd379efded79e9f5a33b05074caf4b",
      x"2132ac00c7bc3a03169585c37b803c34f0031f479327d158e16b0826c607c23e",
      x"3add459756c82b85a93483552c4602d8e591980342ecd499aa321d9a4fc1d673",
      x"fa3805502d9d8acc41247eeae3a354e7c9bdce3278545133ddc7ae05cd9ce5f0",
      x"3d1f0700bbd4b397a5e59bc7ba6e203b94e790358e34bbfb94ad53b6a36ff366",
      x"0140d8a4b3c354bf4ec245205eba6adaaab7e9f2016a0f1f9f533d3a288bbd77",
      x"45a7245b7733ab9357ecbe4a34a56d3c93fa6b172614e2515e9547350c275ba9",
      x"2062b43272e806f7f3ac29313d86243488d0122d6795795f2b8fe6aa2885b45c",
      x"61fdcb8abe091f039a86dbfce06680620716687b5ea87db1b14731961531d5c9",
      x"a6299ca17d58a768d0ca3c6a56b2a8ae2420fcde0c1f8e943bff6bda61ce0d2d",
      x"9a50b60c0d477de74ed2b27fbe4d4196b740512999c881b43eba9181d3bf1ff9",
      x"4d36b55cfd19bcc0e1f15761675fe0caf0a95dd40c735d3dba64e0d919c036e0",
      x"de2a78841ba8c4e095de1df06744fb74bafc23bab975c37212a6471cd27b3020",
      x"86938d198ba55573c6e0ffcb81b228d0801b124345bca3140a1df80d1ff0b485",
      x"a77361cd939294fb17bdc15907e1cb9d6540e4ded71524560b02cd0693625847"
    ),
    (
      x"bf583e81300d0f32d3bae0469bd94cb167db230d47e8f17e994695540031cc69",
      x"33c5fb9dc46f53fd29e17581be5a4390b830f1cacda793de48ef92f225e0c61f",
      x"520d18c49afdc3622d67241db4fb54aafe49f4a8b56c900aa652d50f60656975",
      x"3260ea1ee86acdc475d7141221ef021686e928533b70e156ebf8fb8911560d44",
      x"f73f31ac9833aeb14e79fa4c51e5ef185c85f041dbacd16dd06d40fa5559a4f9",
      x"a130aff85a948c351f0d16640f2ef7fdde4fa1d81a2f79281ca4d3c11da23086",
      x"18e733c1288b33940ea505e400868dd981f9176649b65eb6d5cca1be0e51633b",
      x"25cd46bbc1d595881b0b540dfd636f10ecc19650c9126bb350939f8d85afae9e",
      x"79bef4f703687a1e85f1858760b302ac88767473d2efc90cac643f812e7e28c4",
      x"65e59fe203705db02113616de0e6e555602746aa59cfdc28de156d22c5362d56",
      x"28ca3f4d6b6b9a9d9e0b9968652b61df95bce4bc228f67ef97b577b163317489",
      x"c002ad5834cd01d0e0d66aced04995115075aaea2a2d4d7b09620a1d6171b6d8",
      x"664a58d120dae8655e9d012c3380daa0ed3882aea95fa4937f3676800b158eef",
      x"a425b17962e4ffc16002585eba792ffad6820c1c23f81d8cfaf271af49862911",
      x"92958d72b794d7e4d4c3d038c0948c715ad7d2f478b5c8a1cd19e1bdd9b533b3",
      x"785d7e9bd7a18a83f22cf664c0c9966daa704d90d5123f56a1ce66c3b0030de6",
      x"85162e7ac6dd4af3b8d0af0871262a1c96df37f15443336cd326b42ed28d1614",
      x"c866f504eb666ed6817b7ed1e0d39543d9f92b806d341447ceb01efb6b7bfeac",
      x"1ab166c0f99c07224986e530b4f5feb5f07f6c6017c501562bc87e704b68f9c2",
      x"0bd29fd89c3352fd44f4f7476ada228e643862eac8e9ef5af5ca2ed6d82a8ab4",
      x"ac9165f9f024efd30644ee2537fb01f26f9b979b9176dcab38729a1e05e1de63",
      x"b23865341bc428144148d991fd3813e80b6477a683ae3345065b3bf537903731",
      x"3a8fe20d6b6d0e476f9d58463a4f020006da4a37d1bdf0014bb79368255b3271",
      x"9129df691463a7985fffa863f75575a297cd4d919003bae36b5f589bf325f71c",
      x"79ce7d72011e83d898e746af2c509b44cb0f7963c1f0e6360b435dedc56350d3",
      x"9007ad57096ea21c36f582761a927d0cdce7a0c584a52d722e7408e0465f3e76",
      x"9f59b1f3a43b5b2e1ae3455f77dc4f06c54d45d48e6f7e4eba0eeb27a492c0ce",
      x"f659217140ee5fbaa7ccaaf7f9fabf2c260762e5095fa1af846d584b7a867914",
      x"eafa0f430c88ab294d7e375fe47b249b89a7d6efc42accf5cd02091ee6e13450",
      x"d8fdabfa5d3c700eae00d58f0930cff26c8d8802c9416ff05b25004be6adc216",
      x"6f9889d3351483e0e60bb6d103570445b996299a8d79e20d8e30fb6e6d942ef7",
      x"20c59db0b339ccf573563c64eb09f8d270d3f7704482c9cb6cf31c2bb5ccd558",
      x"1f9f094560f4302edbca2879fa4d39d4f8c09229000d84de8e8fa6e814d36b87",
      x"cc58236f50059d3e21833563c133deab908b1a7a361b76656619186e8307e453",
      x"bde616869d48af66d61b3589d11cbc015f8c3ab10e4f6246e05b80308cd5a936",
      x"11472df06a50594f1e17b0ae5380167d3f6b7dcd3049b5d940172064dc8ec593",
      x"d47b923d121a25c54d627a5d6c19b5ddad2c9fbd8e4c35a1d89d3dc492d9ad01",
      x"1dfd96d6f7a3f90aa790c12e9951711b34eb43fbdd9a407d30978cd614f0a210",
      x"215e55618f61f2268880e01d8e40a4fae153ad273f145745cfb8ef1fc38879ef",
      x"54daf6932cb8b8088ddf9c0817e65707da1278ccac92170ec564cde2dc0f3f1a",
      x"18fb334e0fd628272d37ebd8205d6911bedbb84c8af1c6e5804d766170acb6f4",
      x"b33a978b205a2008f67b30e33ec78db933c29d094581bda2108157fa1ba9678c",
      x"4a84d8015db40560a7a921e5a28a4f17f6232d5a666f22baa427ef4290cd8b54",
      x"18a00a45f6ecd28cd9dea64e5d85916fd05a9788c140fc5920a97c3102a51ec6",
      x"96ac5e7d9b1a1aa73a6e2e99e66996dd466e296d81dd00aae20157cc14860948",
      x"ef70f59280466ac875001f264853116445b37cdc678a52c8a2e39551a32381f8",
      x"dbfe29e59312d6fc5ee790b0ee7c6e82d59e624e04f90cea212b00a506883296",
      x"805850c64498d9adfb38e67b92cc7ed8ed4e570b60f3bf7415d444fb397e1d0b",
      x"15de5293e889ddd32f6bb54ef1cf258e91730ad6a348df97d23746fec05d99ee",
      x"317c0640512639eb14f9c0615fce7a38419772469d986be7d9dd0925335db593",
      x"ebf239ce822205b25a6c373d85f27ac21d155d7de7386e4de9af3bc5438c2dc1",
      x"9be97799f9bc5185416acf9082cbd4985daf030dad66cb34c50a2335c566953b",
      x"b7fd897b7a58395b2f0d9fe3f1dc8da3e92fcfbff8edb73d97e41e4001b006f8",
      x"d2eab40abdbbf9c41b1f6c9df214a2b81e434baf404506a88cea5eb2beca63c7",
      x"8a189572ebc7e9ed0b23a30e289d549733f5d4a0466f45c40dbfade950bc8be7",
      x"63a6e48f45376e15e5824c95a24886f80e77d542b9620bf23855d8f0f95bd421",
      x"af60486e8d2fb4e050326acc89c9b64810a68eafcfa855e143128b87107ec1b4",
      x"a39b389e7d29a0dae055efde8df31d6fdefc34e49c8ecb86726675fa6bc56104",
      x"24b8e2dcd98467f0648039e6c9baf1f58089c100ac4260775a39ede40be99da3",
      x"36394df3e77e688f9d5a157fe3289d91b88962900e9379a9eda9c7511e9b47a3",
      x"1664a8b746548e0d7838d0bdf6f5a1b111ad76dee7700bf9d24e1701fcd863d4",
      x"db5c455f954ff73db2c44bcbccce60a7b6bedf8fe5a7d80a9d57f6efbab906ed",
      x"6ad26f417856f39c66fb61c4d594506c9e03c087630ed485be12ed377001e379",
      x"ecb8e9ea979ed750dcc709915acb0d9c9c3e6d5315367f662e616779f60fde7a",
      x"a737dcbf55c7896cacc1b2191c0aca23bcf3768bf69467d11d01928fcbc91359",
      x"d53bb68f41eb2ac2ca5962cda41d1fa04ad172befaa8a3305bff4943d477e09c",
      x"d9fa7784efffaf38de5db00a031d460f0af0703d34a35817a2a4654271ab3003",
      x"4d7fbe303491425888853f5fc1c857f966b998e6396c00f77686ea9253f2e35c",
      x"fcea357b3569420fe65f7ea2ad77013f176db4700a2690ce468dc3a1fb903911",
      x"22a50832a6a8b2be8125c7e92f2fc1d3b98d87d2df201ebfa93b591997ee2b6d",
      x"82741b0228557e518bfbba3aadeef55a684b3a30dbd3906dfb15dd89e1b687d1",
      x"7526d1736bb1e0299de2aca1272d53d436da7e88c6d892c21a3db52e4a56a33e",
      x"ef5be9a93a4a774de2a0f084dbb54d1cc58fe2d3b39387d9c75bcd89fbd829e6",
      x"7858058060b8334320c3883c6a88dd58e79b29068c7d18610d683fd80c478a07",
      x"8cd24e5594764011e45f41db74e9f7397cf1add36fdda3310c3c33b97c51cb26",
      x"5c40d258ad499b031fa84af6e5783d9424cfa912d8141aaaa52b69115c0eaa90",
      x"04ccceab4e18df651016978d4b9d0fa6b05f143444ba74f97edef6d1e4c82d17",
      x"9e013f70e8599517bee110ecb110c777bb6f893280f6aa3d1acdc7ce8fbba4bc",
      x"80a20012744c5878d1c7c33c955256d172158ec704e24f23367e0796d734b4d9",
      x"ad1919ad7e63abce10c3a634e000e09e061e1b2f969fa85e6007954545b3f0a5",
      x"da7a5a15f3f9b24ed9002c5cd3df08b1b8d1095f367b471cced339f3ae570f14",
      x"81b290f4a618a2998851223b574a0d9640df44b241e48cd35d8e20fce1f55bb1",
      x"90d4087847b64b802f78ca8edb3ff81111ae69d5658f0ed2ccec553d8c2072a3",
      x"5b023d4ae988993786c65390a70eb389565d0aefa8a4b107712bc9de7c51927a",
      x"116e36fd0420ccc5307c188e5d7eabc28f96c6ab8c77a6d3af102a0d5df7dcb9",
      x"42fe2808989830d69119f98e4cbfae14304a5137ed0e19f6c9c37ac2851e67d4",
      x"0be09566714c72d57101205b1f1292f2211bbf65786d9b1c574d5d4473930e2d",
      x"53398f954a8efa4e6ad96815e92372505c0a25d20e9072d7fc880ba0e49ccc0f",
      x"37d8789c6a2850a76b4d4dff93dcd830041ea9efc6ce0a1fdc3813b0746b8b18",
      x"013c1391d138624d045379f3a8358c9571f13560f09d9448d657002dd206a7b6",
      x"9f06cb64e02d1f86c68af0bd6a84d4f651c9ffde0b7c17d42572423bb7e54364",
      x"12b250d3a13cb04c3b5c99be761ec4aa131c64313f6a93246e39a558b09baddf",
      x"291d44df5bbde98caab6d825440cf67ca3b331b3297beb9400bab9747c47d93b",
      x"16dfb8331dfdf7e92507dce2c1e6927c396f6411dc6fa799fef17d45d5c3e85b",
      x"464b00269cc5373089f7676d7d16ff786b4f97af7fbcc12748fcc5fb619e7ea4",
      x"8507dd36bd681a3b9481dcbdbf6ce0528636c548c77f4230fce85a4f10d5c4f6",
      x"356984f092596f9c1e4f92c59b4a121a7b818cd051f4467ac96f10d6f86af4c7",
      x"86131d2e79ecabd1443b8210131ac155d8079a49f65db8c92f2e53b509734dea",
      x"8e0e92e485a8de09002be8607d6f95eb435ce598b348dfc116be27f1d825bab1",
      x"6473041834aa1280feedb59a6c845e2aac254595e441e62d7538ec2d0613c874",
      x"4e8c7f22812ddd8f051fe597458a122b0005efb701fba7e80d13bb9fb1bbcab4",
      x"c0c3d7f66718739999495c85e2084f7dd3585b8972c829f27d95a38ccaec132a",
      x"6a9510f25197a9d200d45cee5671a0263febe8615551acaecaafd8153ddab909",
      x"a0e7ceadccf7b15a557712e20614ec8df3b1a74c923044f2a35b49bad5a3eec6",
      x"f113417bdc7fc0ba6115bc4fee0e9784950e79b268e5148a58104f2c5771a538",
      x"1611cac8000b86f98e70a4b11614bdf1ed95894bd69e81bdc797f45dd503d590",
      x"b216e59f7fbb134b4b1a48ec1bcd5401942434c495f882a53749eb6196372840",
      x"7ac162dc63436620aa7d941565148074e7aed6baa886fcf76e1aef7761a1a00a",
      x"d555aa70ab589f3f407b86dfbbee3c6d6d691c77749015b47c18d3669c6a31fe",
      x"c233534bb1c743eb589a62b63a953b7faf7f99f615a72cb215a26aaea2a9ed6d",
      x"c7b78f145777ae359e871258cba67823c7d3a25b2dde78c06a64bdebe9158495",
      x"4ab7eb4c89e95118fa8874bd0ee59aab264a87b9b1c0138f53e2f6af222c8504",
      x"afa5e380951c5740195468962bbbc6324b34b610803cf126c37480f64e5d30a5",
      x"dc2325d0abec88d95d872a6331c6823d76b7b40a309985f2ac3efa570b728978",
      x"8cae43081638367b95af2d9c0ca8972522a7264a9202bfdb7be21b7feed3da86",
      x"01523086fdc6c1101dd0f10a25ca2b01fe707580c9071ede21b78117a27bcba6",
      x"cdc2715cada1ae8f622ff2b870dc24fb7f70bd74831bed7db640d5a2ca7a3984",
      x"ba93fcbe2f63e5d41bfd2dce9373255d091db5492dd1d50ab75bf5d3e1848f02",
      x"bd54ee0e99fcb82e322c5b547cc9400c7758863d2c56ca2bb53392cce26b6639",
      x"23ea363437ae47ea873c3b2736fc88d3ec46b53c0d9216e1d6c7fa7c619ed08c",
      x"18ae6167f004c4a0a78be71e169a512c313685f529c22e09b038c51300f84b88",
      x"b3a3a9ce68427731b66a3148dfb8c0f2c9b9128ad006c325db3b0636b2abc503",
      x"eb9a738a31d300b8b06f26f16cbf730bbea37eecd33e472d5bc3860d87ea0212",
      x"d0772438044d1c5b7d58685f8d1abc1feb72a902e16ecaf2f758809cf0c22a6c",
      x"156038fe4d494a8b80c2a27fae3392626e124775f99398760820cff1c76de210",
      x"bd8caf6a82232e932f9a1f8ccb6c80bbf673fe3d8ebf595a6ae79653551c6ea4",
      x"ccc7928bfcc0477d71d56d6f716c66a1efc8d11438d3b75e15cc7e61a062ed1b",
      x"4ad604b3239b750b1e2968da59020c0da69d47fca4a377c8dbfffd8eb0029a4c",
      x"9c2302d20e12095cd9aa760601244f141883f5f4a48f80849be18dcf469a3d60",
      x"37ce666d9c59b8742e77ad6e2ba230d87c8996fac517b5252673047aaab5ff27",
      x"e85fa5da2dc02aa535e78bf97043fcd9b5fb6d1b5c43b0571ab819b0d49d0032",
      x"21e7b557b99b8e5d58286b00f4b41930f43812d9fa18a3daae4e26018529adcf",
      x"d8038668ed3cef4fcaa4b4c50311323a27a3b9aa0c388cff6b6650cf5b9019ab",
      x"a5cd177cb19316a2e342782d206841061140872fc5210da9906e28fef8f570e3",
      x"869d0a37e4c51bed00bf1633419967353920ddf7e0dd1d2989bcadfe6f345ad3",
      x"e17c1ac790a4f74ab1bf322f20bc81fd87e6cb77412cf214b9286464c75290d0",
      x"9c83d455a7e41f16c8b1af89515d5ddb27e67d44b2a2a3ba32425131cec71289",
      x"6064ef3c9a6b5c34d7b334138ab7b3359c4ec136c159ae610d1a5d7275bfebbf",
      x"8e136298ad4cd9e164755ce0813e448416444c082cbe2f779da8a1452e5c08a7",
      x"9c8ba2c690f48355cd2960b2b2c240fa4a867e74f667262a221063446183fafb",
      x"3eecfd4ba6c04947657106ce3ec404fb7da5e5ecfdf917a168ad91c806394db5",
      x"bec97f3cec576ac96e0e4891ffc03aeac5a68d6ff877bfa02692299ac89f0643",
      x"4b1b3dd208628bcbd7f4c01e4e4d75e40c7d16e2faaa31eac7230fea951f35bc",
      x"8d9a2877afa0c847f441747759e3c58e7e5f0db07ff4ad2d70409c50f5c73226",
      x"4766ab08302931ecf170708aad86ae5d5a1b1ac4e943ca9a328077f127dc951b",
      x"2536228ee9d8eb252281fc146e20c9870988320a4b680ff24fb49b01e55c690f",
      x"1f2bf715d7cb7c6258828b0902fc5fa3491c0cd30109e8a545f2e477fb8e85b0",
      x"d6af4250216e0b24a8932651afd229f0aacb4dc6dc7011fbf90be6901f214977",
      x"94f23492ea60338bd9feaedba7bf6af48f1b0c90272f69e8c08d191d5c7b30b9",
      x"6f236f9212696746473d02cbefdd17a7e1d930c65ed331c65b5d29e5e56a3208",
      x"f0dac4c210cf28edda0a9adeb5e9fe5e1e657e94da910b497788e629b3b5a689",
      x"529912b4c9561d61df67265bcc2314d84efcb4de0e6e206153e20a874edee43d",
      x"27dcf41ee6a97b1bf227bbbf140e9624d08e314a816e4c948af1fcf0d56d4176",
      x"c6f1c81c0afe6cf1a7129cad72b8677054bbeefce4ec51345bf8c984f6777733",
      x"340cf2e19dfaca8dd3521ee190311264d941b9741feac18f7d297e7fea38419a",
      x"f00a5118dba40dfad2c3c01814c18decc98abc5343ca5bd5096d8ec822ffd772",
      x"cfa3bf5c5a6e2fe5b57949b138e8c3f8f8d82e1973c55d7462820d7afe0adf38",
      x"92955c5fee5965b3073ecd5e3db87c0880f562f785b56cd476b35d27573bc4e6",
      x"81ac7a6e8c90d8de5abfab61c357baa83ccfd7c8a6d188f24a705f0954ca905b",
      x"b49f70bb8e8ad9e4f66368813a70bb2b574f941146155da2a864f8ea9c416868",
      x"df5cef457105d52fd02bfe73a201b71168a2563e7a2153abc0d417c72342ade8",
      x"d1dbd088a94b4ee06d37e24fe423116d4cee52753a74a154f0fd5b8d67bb96fb",
      x"11fc7c3510eb80161565878dff0a3c0195c5c24a066d3e02fffb0174c0ababa0",
      x"5eaf66f65f8a1863a4f500cfeaf708ad3609368ceb4b47081f6ca7bcd8b7b5c1",
      x"a9334df49348be34e58fbdfd8a8ef0e5a08a715146126f4d447c0835bfd5c0db",
      x"041b5e835a2d1292e71747651aa59125eb22da60ee7da3e9f4bfebb933230239",
      x"11c7a4cd1ae6eda7dceed9124809ad1cf079b24ef515b664b5fe6dd57986637b",
      x"a4aee105438321be778ae144e4550cec420d39f65c6549bc627a5cfd7a5b52bb",
      x"c2d5d14371cbf0d6374e7ce6191d8ac542d409f8c4d4f81445456457c8c57eaf",
      x"8b852b3a589f7741fb424a1ce54c5f4b4e7c40dc07a4ee6e8d7b9b599c7cdee0",
      x"13f5d6fe6dcbd3cf2512989a9f2e6a41c3ca364cdac117e181df6e67bf6e9fed",
      x"51693d01fbc21a3364ae3d20700ef189cd40fc89382fc1ff8c073b2b47e5a6a0",
      x"2045fef4d507b857ecdc2b439cfe07870042e0fc4f25cf94611644f6d6c18933",
      x"883d4aef1f1e40aa04b6ebc77aa7b6a168776ac0708a9606ccfa2e6e596a2564",
      x"35f7c96dee2afe549de534416d00faa3591a873713ffd1e2eec0e04feb2aa9b2",
      x"2b5d8f2fd3cfc6782e9b0986c011c4c225873af1b8d9e6fc9b79dab323c48984",
      x"163b1d000cc293bcaa2adbdb195b789362ac58e1b621cd6694ba862a53bdc007",
      x"5b9e3122b1315ffbc3f4f7e2303d095b71f42e85bba69a4f2cfbb17fcb39cd86",
      x"2ab620c19deff6fa8072705365199b5f3f07a841448211290d2c89f509458cfd",
      x"5098e91c9649514a6bc9206e2778bf8240b8be5c5103a0bafb22e41df6c8e1d2",
      x"9d8aa515f3eeafd94c02b9caf42a345959d6a2b728cbd9b0ed6f38f79dde0326",
      x"f0558867e4817359be72ac85d8aa52730bd8148b61445c21782e857b3acd65a2",
      x"6a1bd54beb5c4c8016a44a5ef56314a834551329f9aae08dcee7bfa69530ccc8",
      x"de2554e6b533c4d1f7cc12a4a41da29674b733332dea7947d98bca641383befb",
      x"b260c35ee7febf672cb2988cb606505e22857e1a6b20382fd1d293465eb9f084",
      x"1fea271e177cbca3439a6b027c7bcb7d81cfa8d4097c0fc5117b6eb550431a2b",
      x"12fb6f39c197b44667e59e1f13c30615e2013e5e135c6038cb47ddeb78c71d59",
      x"27a13b62accbd708a92fc082c7b667486d7d41c850e0acc12cbe4fcc364da560",
      x"b8a208c147261642a383a9311c1a2dfa6a8450d27d092a7df2500b3b0ac0e18c",
      x"d63c023b43614f03dd521aceec63994538a53c9138d7696c65993ccfd4f556ed",
      x"895957ee2893623fe4a58f38a107ba0947b9a308e06834d51027d5467e099f33",
      x"3c0fe7182053ae0d4184fa7311ea3791c769bc866c44a4abc92be376a36a5185",
      x"d4f26dcea8756ce194182e2326e5582cfa385c27fa94281887b07099a3a6e14b",
      x"d83de44294110d72d15257767b279553024dcd7bd89c6db723b4b7ed3a15ce49",
      x"00cc6b7d95a4f9b028145e59e07da192bf59ebdad588a5bfdb6f3c390641ff5b",
      x"9c42eeb05f3b362f1fccd5fc6c08eb4df4056a0d0d146141fbc35fec7123bf6b",
      x"d06d3bdf533dad8d7a8ac30eaac95373039b8f8c1c3c5a681a07cfc3b23f929f",
      x"0308b208788395471b030042d0ef95f7457fe2be942c2ba0c57763ee76badc51",
      x"81f8b9966685a987e1241f913e3206188d6af8a256e761bf8050627012457c03",
      x"3439a1ee7533ad0d8675f4c26420cfb7f08469c548a06e47a6208c589761f28c",
      x"3550bdbe8b86daec83b0799013694e0270d4e1994bcfad8a2cb5c7b1393f9d30",
      x"4869a7288009de24b69e58cd1e817489c9de545c3cf7d7f7effd378d39fd26f8",
      x"d10034a7d7bcf5701fdcf9947cdc2d6d9fd864cb6d7167684ee4cdd6d51d1f4c",
      x"6bea5a3ae8565d51611fb1b2b6f16a3d7fe20fcef789a02ed869f1d3138c0767",
      x"231931b9d3d45bb0d59f22316f26cf9308fc349c6b698441cc5d8304392197f5",
      x"618ccfd10def017ae040e953a2c04294ad95c616f674ed0d9969bfa23a881884",
      x"944f29e33806865d3c8c3e3920ed5b498035518b39a207e640e7f62ce74c6262",
      x"0c64bc66c2b0caaaba1685493b31f0d249c6a1b7c3028c729a852c92f54a25b6",
      x"42c877e6f40d915a962d449ce409f74199ab964099f5f1000bf347b0cb80d930",
      x"e36b4d88c438d3bb277c10a546664bf6d661234fc56f604b7a484d481c505233",
      x"d0cf9925e4b3131ce2cb136585e3bca9b662dd93fbb22240bd383605f04ee72b",
      x"f18d2a479ae3e20ef7dccac0c7f326194d23732d3249cdd42b8eefde7db0c156",
      x"242c5c2449a79cdb3003dda72382f654003f8899ba5d63782fc2d2c88971ec03",
      x"195ca99a8718e2b0eddcaa5e97d9e82757a58cc79b9bc9a69342757b2cfb0f34",
      x"d8efb0482fdd7021ce886373ee6f3719c603bb373eadc7710ee85b8622b2dca8",
      x"be1ae0b5bc77a2fbf48cbc1230a902d356744242c3b6ec9b871cf0516fd9a055",
      x"6c80321c989555a19a1479e94d2edf95a417682c0130524a5c5a65a5957d370a",
      x"05df8c39d15eecfdbd566405d6622cdba80cb1179f281d0e87bb24dff02ed02c",
      x"36f5cf829deb309777f85de880f009ec44a866b4ba8be6a7663b2a2f9dec55d4",
      x"a19945c28041f9ac542d13d039327d6d72dd720d3acbc27da24f436dfc54dce1",
      x"a1c08eda443cb06cf21c0a57f9d480a0605346ea3bdda660bee06c2e51f5d27c",
      x"cfaabee52ce19a646dc7a38910973c4b78aa2a1ce65bb3e8b5e9a1f104bd11ed",
      x"2cf3b328628f99bdf6c75557114361c591edefabc497f42da41b23c1624644ca",
      x"4db76f21fa7dfa70fa556d4b639c6d10142badabbc6b64e4f1f4c027d33e77a0",
      x"c2aea497e7f8647390f249c3115a64ab7549bc3009ee4a8353dc7983b641228c",
      x"d7df4fdbb34f71350d20437866109f0ce3d88d4ff35253311cb8c8d897c9d966",
      x"1d702203e76c786d9a60c21c34a7575e8a8ee58e57fa540d32558707eac077c5",
      x"661a94c071601f7d83f44504b1a5a8ab9fce43f4f038f012e14e09a76f5d8f32",
      x"6c94c65ebba894d2dae64ac4b64e0b4d2d8d03a6dea3a8a905eea917364772d6",
      x"0478f8d7904d8d5d23905d77b4eaa1896180b1971aac67469783f9f8560125f2",
      x"f968d91b0f858ef241da24b1e0e34a80860818719579e1ed22500f2750e06eb5",
      x"9ce3a2745207ac7f41e8d78b8f23994de68c348a0f8b7ef448e2f7cee9ad6494",
      x"775d514e5c254a41a014aeef6dd07ef2dc6de625dff7f6c36622f721d7afd276",
      x"bb7aa4a5d5153690c7f8247fa9380abc9e43bf541bd4f7d00af2265ac1db7661",
      x"a4cdd8f28a2ba1395b8f20e3ba4ec68670cd978189ffd4d099023beb7690d476",
      x"4a62901c46b581ff83d02aca58bb664c4ce69f219dc680959493611261af389f",
      x"b1177894c7279d5db8e8df7fa0c9debd30a4c95d302792aa3439b70b3b8a27c5",
      x"1c2561e86c8d523c063209dbbd1760c942e633eeab0abee4631526840a48f9cd",
      x"4abd06899d87d14f90e1306b25057440720c70b62a366f81bd14f05cee7d355d",
      x"0d197da4f5dd04a505d0253a2c5e2194c1b9877acaf54da95bad52bd5d0f1f70",
      x"a1227d2f1f678bcc8c30584064252b5e07f385bf73b23e1122df60ed19977d5e",
      x"d40d634c9604c645bba6f3b7a1b28772f10f245a511b3b51de045c657801f3f1",
      x"3e21d341e9d8249cad573f95b11914af59e460e856442e6e1723302a904d3f28",
      x"57ecdadde7c7d77cf9c53738ad531ad60fb52ced17dc45420a5f4994f75c90ea",
      x"f716ec676ded6580febd2dd1777ae04fa165719d7692170df3831963e8c68dfb",
      x"448128209a6899c862a30516cd88809ec14215f9d4f634090ab69b7e41cb297e",
      x"1be9bc3db7e0f8c4430de9c3a60602dd574f4d6687851e9f23ba4d397c72d82d",
      x"05dc866e8f8e7f7c7f37949199705fe4b1e393c4d4e5d8003d3a75724fbac9d7",
      x"d74b7c4e9fd657f2eea632ebc6c44649b2c7d6a734db883a8b42c1506c70d8d5",
      x"05d2ef76ac16d6f022f81a63093f64a3b1a307756493500b788f0ed69af0a3eb",
      x"85200445d3eaef6e84a3893be7d31f2b1f25a967f009821748b9a2bd3538e0b7",
      x"e23f82732ca4b6bc5e317a979e7e00e1651ef93a4248305208473825e8d5b973",
      x"461e4a982ce69418e7d6eaab768e73548aca78cbff6e6d489d1f85879f0135e2",
      x"1107e349140993b864e58a3bedb750b6abd8ddc7d43455c3219dda246c8355b6",
      x"eb68d3806a1c207e218caceeacb6dd2819cf0c52bfc9db6367fba8e9fe1a899e",
      x"e26339be0827830c74267fa730edaff83097ba74b5d70e5aedc96d828ee23cb8"
    ),
    (
      x"8eb5f9dda78774385ebc8a22d883c5feb2f6c7c01b8ccef3e4c886b44d079b68",
      x"fb8432ae82a2e3f0f83292590eb3f1908a58e974f65905e77892ad81bbc955b6",
      x"6fe00282aea2e7bf908839121ddffe30409c70550b833e2c8c986ce416c6f166",
      x"bbe98643f9782e2dad358ff2586299fb3dca05cab2dcc4bf40123ac47a571eaa",
      x"30be63aadd5281d96c17e247e2ce719073b60c0d9631adcfebf7fc41da8e771c",
      x"82c6abb4e384056f98348aa7a5b863dd08b58988c1bd85eabe784cf82f07677d",
      x"8677064d65cba2eb132ff833a435232487f47bcb2a5ca0b17fc8281169db0aff",
      x"51c457e7ac11b0927a6875e7e8985284e1926dd2fa62bc07470c6938d09177bf",
      x"30bd0a3ba7e1548536d93aba2179654347d29b0b01b6d127dde0726806472a28",
      x"c7c16c00c9b7ed94432278adc15eacd95ad6f3af903d3753c54a6375299dbf7e",
      x"fce5fbd5729c894499883bf4ac3b0a65c99ed3ca2ab73f7d20fa101c031867f5",
      x"61c72662742009d973c759877e10a85b9e8449a4f53edac5e8983d0f7fefc6aa",
      x"4d515b65b12fdc8efefaeab449c476fb6555dec5a51b59f132ca34972707b0d7",
      x"3fcebc9dfbee2c6745c19af84f9131ea6472201c01d623c35a90c46175934428",
      x"aea968a28b7b162813a4c142a7568521e3cce7d8ba673107ab0af1b6c2db75ae",
      x"71c0d99a825fc72e5931659281cc4ab6bde44601eb29706dba3c3fc315cf2165",
      x"8925ee26bde03d48c653fe5e903e64465ca2f858805a58db7c4df021335a6c46",
      x"4a2b28fd7e478d3bf179b81a1e215e6f937866ae25810c3a761b8b17d030d0dc",
      x"c90325b8f48982a94cd0097f667cad27d787ada5e95cef8353f74a27ec22fabb",
      x"2fd7a78af87ecb574e0b8709c144679bb215873d1e1b76b00400bc1223b92663",
      x"93c67374f0d8ebbdb7f21f1575992ffdf02cf9b6cfe10726a9b13f490a555c8c",
      x"c39d992a33ce1670ae0f6a92bf892a26d15864df1afe90a47aeb489e4afebeac",
      x"dc16a6b29d44e4df9a8b9e076890a5681189f9f935b978363ca2a678495fd335",
      x"474495ebdf20f9804405fd468b7395cb97c5713c1b10c398acc8e94e28d780b3",
      x"18eab6a068c06c0a47e1075c7a5e6cb33ee48c6bbcec54a2e8d87c3b2bd13bb9",
      x"a78472cd9e64c4198b77b51104d7456e206fe48e19276d517623df880f71d889",
      x"31c760b43a0216ee37d42d880608d4179b395335c2d71467a6b0dc6b0c959a30",
      x"bb30415563ae1112ef862041e978675113acf5b29d426aff888f0a49ee02600c",
      x"33d3facc7fb95c0345301d1cfc9d6f1d16958d8f15ad62c35f68278251c2d187",
      x"beb081669aa0a5029891217d1faabbe871d2301f54dde1759604a06c65674f26",
      x"a4fae5602d9183681b0779a75b40cb23249c1aaef729fff2747f2bebf51ce0ce",
      x"66ef969be1e472ca1b5fca426d69ddcf70520086d78ee0d6f7729473781c57b3",
      x"07255217d8202f4e8ec44af6b17b7e0f021aca5959e6c4a994e0dd8393796c20",
      x"eb1256ebab7ce7238247fd60274b9bb871828be74ceaecdf0d885e82351f7d52",
      x"2ef5b894e10365f4cb9d7a67c26d8676d20b767227ceb2232b466cc30feff0bd",
      x"da030b6e038d5f40e40e2e429d48d7c3a5557ba8ff983ba62f178d9d04da4d63",
      x"bcfac35a19d27b9cba5e974692b583880bced8a73ec86a924e740a6693bc69d0",
      x"15cc9a0fc20959690ac78ede8a2610a08e2859403f226e0e82dd33753dcb3eef",
      x"5f42dc8199a47be349c91c81b1dcbae95295b5885501bf1a028b059d5514e87e",
      x"dd83de78746bfca55999310c1e837c7bea8925327b47351322df53316075a142",
      x"352e83128956caa63302963c4ea808bc3ddfbfda55cb413e6e2b16866a9fc72b",
      x"4677753de011020e7de3f93ebfc5b5acbfda5280057641b65aca17ed54a879c6",
      x"365c40b59bd1c38098b14f0a4aa67610cf35f31db34868884b35acce42e31a14",
      x"48686c30a168d685037f44194474e9e9ad618b620810a67875879179ecd4faa2",
      x"fb0a22a60d63c03a460c82c4b018e500f2c6509c2cf0dff83e57ee5e00f8c067",
      x"097f50aedacc905280056ba8cfe2ee44c01becc477001948074baa961690518e",
      x"ccd20061c6461efe252c4c31682b727f35f8f90e59fe869dabe59fbe1dc3b17f",
      x"cee298c995fd5f5b0c5fd0838522308aa2075ac33f835c5684253bfa08738dcf",
      x"07444110d9b6df79f0c91d6ba394aad111a3a31d331101583aa3a5dfdf74cdda",
      x"df18a6bb27cfaf6965252360fad0ca3cea997ea31711a78a642c7ec102bcd6e4",
      x"3dd6a9c528885eaecf2630900c43592d7a467fad5eb267435123f2d295a1bc52",
      x"5251015f3e45ac8a65cae1fcfd53e54e734abfef4ac9cdd127fb524f5c1dead3",
      x"e491d6a40665a59920522bad2b92c393505d381be6097a8fcd42f99f4f8ccef3",
      x"3036b9d0fc3013a56272b6dfe796e2793a6dd68f715cee99c0634a24f59c7b95",
      x"134b95865e1b2697eb49541ebcbc0bc7ff8ddcc8b102c734d29bba49add2e9c8",
      x"660b153b82c48061761294e1ac47ecc2f95a050694bd9f4ae0859be1f6b0373e",
      x"495dd0e09bf8386d26480e9d51cdec930155b3756eeda1dbc6d91fb6346cc692",
      x"d24e1901234d4e5aa8e601393f5f67f16bcf05b87cbfd05bffdab1b75f5f15af",
      x"83318250a573a3dc3fdcd56193e1584069ef11ee77f862361b5362544990e6f7",
      x"42eadd03f6825a0a8b9b4680b2add08a1a3d58810f9f97043e9b6447f8674e97",
      x"0366466f21501d871d98a5dcd6f8dbb86fc587dd257bbb9aab68931f94cf5d4f",
      x"08a4480d64609ea825833c3bcb72b5a65d38e31181095f317afdb04de4193252",
      x"410e16543de953fd60677456f1834036e4c39df93deb4a64f2e2c73cedc731c4",
      x"04a76560dd1af8d698827674cbf131a369fe2404f378fd2b924da5d73eb371ae",
      x"130b7b0a895f5d55ed0cc2ab09343b22d9204a6c52296af2af714350b481108e",
      x"df282c0e4bef9b9310b229f9d908531a4286aee403af0570ddce2b242d2ecf2b",
      x"e0eed8ebfe47ab311bfe955fe3851ddf9b88f90fda6dc754ad5a2aa65e9ac1a2",
      x"c2346b5740a125585ea76af2e5b760f9c197425c00065cf6531abeb88a8a6aa4",
      x"358e0ba22a6c6f005128adf449361ca91a69cc8209c1bbae4c5122acda91b572",
      x"04ff4c74aafc31b603c5a969d22009c742d0b6f96a12b2cb4e0eaa43cb01cc58",
      x"a49a096e9c77305312c0cec277c2dbfacb380238ca1e3795771ed8d8ee24d378",
      x"5b8026c6aee3f38453c104bfbcaff82ca50cb06a20eeb23e0e55fd3b13769493",
      x"320a55dc6559cbf39c207a8d8cb3c24fdf1a8fa1b857c66d2770719c436f1644",
      x"0d015034f3c25263309eeef278a9caea607f35d3400f75551a791231896d73c7",
      x"db349af6514ad34aced46536e1853706ffa0ae9ff7ede6431a5f35c9b5778529",
      x"4c848a8a04eeb544d8e2825d7dd6b2c47f15a1101f1e248a9fdbe29fa306a836",
      x"8499eb0a4a5c9b165e75b67f5700872ba76e8b04a729a6f4ea0b49cee78ee414",
      x"5068d559b3b12ea472370d1e76488f9bcb36c03ff15441bafe94a5cf20db9cd8",
      x"ed05e58a3ad9e297e86f939d4cc87f92952d3da2e7227cd8083b468ab739df45",
      x"0073c58f66d6712a7ebbeb58125b66a3eea1a507a702108cf15618a7787fa27a",
      x"544515d9c2b2bf949f99cab281ef57fe61e3ffe1b6038a4521c418c82c52ed4e",
      x"188fbd32abe21bb7b09214f68c995c463fb274dd4215c1d679ef39125f82169b",
      x"e35529e00d2e3a07510b8a2e3c95e1d32889a0f8cba720d93207197d06f15033",
      x"2de91feb77895d71899b2343b253e3712a05871bbf05d2efcf86f28505cc7d5c",
      x"5cb7c2b0a90707903a7040075d803dee885088e42e5b31f4ffdb7429c1e2c638",
      x"85d49b15e5e6b74d923c912788b279c89bb9be1383f8711bfb4e50d260aa4486",
      x"a74b9af7e698aa27c8b4800466fd9e7f694a86f07ddfc9becd080b3bc139da71",
      x"87e5f53b9cbffaa356a7d768664c8327081f9bee14482e02bdc97ce0f14e6ed7",
      x"9e01f74bc6a17d8f85a7777c032409aa46eedc38b5898740328926c681d55dc1",
      x"92ffb57ad546882b34b4f40e76611d1d6270c3f362f2eb774e318583a375c078",
      x"440643626527b9ca0a297a1b5d4ca834dd64c060de9aceb1f99ae5cf21759049",
      x"5a61a4485dffb4a6336bd17d2e43abfd70b482bc5876e816100858c1b0c8f14b",
      x"cbbba3eb5e758342046696b71a06c43d7119e8773f80bcf70dc27ef5993a18ab",
      x"09694125adb1677f61b92a4943d3d941fa669d36c6887148c3f848c702584614",
      x"7070a4962cfce34e323732963ec5e6158475df11c19ab2170cc50e33653f8d2a",
      x"4a96273300b19ed1ae61b61386833c74282f2edfcfac0f39d5a9ac244564198a",
      x"6d3f399b7436022d3f9f6df3a33f8c72a46cf7b35bbf1edf44468807fcb198e8",
      x"365fe16341259c3045666d44df342fade0951712d90e4cb648a6c4fec4a0105c",
      x"68d4ac362bf86b8e22db9b122b4887bc68e3b3184dc4ed75ef9532eaf8ea94ce",
      x"4e650defb361043d79953fd312fdb4de809feda0c828f435fe922463adccac6c",
      x"87f89fc7ac56ec5dc96ce95b31fc7c60838e6ac37253076fd860a066e7e02a74",
      x"d56fae5bfa9915a05a0a200e9879ba4322b4f2036135c68e1389f7fb0d24b0b7",
      x"b369e8b0effec61b574af00493a2df45718fdb08e5622038fcba3a1ecab28e54",
      x"f52b97fc9ed788fe8f018591b2d783c19e390aadb46db2179a92a5d73a246b06",
      x"6435a6557bbad66c667f7a55e196aed4739534ba6068e9e538285d640a692ee9",
      x"6dd99ed35c7442ccba55407d924a3c2f8ead481afb902f6a160cd0917a83a86f",
      x"471e0db07ce6fa50f2cffd3b457681e7cd6514760c5f6654aced5435ea2c1c25",
      x"09aeb8e239de7515a1a3cd47722099fcfd227d8ea6cd88cec6a213108f25bfdf",
      x"c41fc4fbad7fa70668f6b5321fd543c13613f950cb3fd07d0d8fd2b1b544a25d",
      x"e80c9640d84a6580cfcc4c198f5d644c6b39ff9d6dcb8cf5e2d7c83b18fbaf33",
      x"8de3cab941cae3d3efe4a1d4de2a14a3a0845dea4d6012e6a92507c5461195d2",
      x"0ab0d57299a6a4e85c391d4f2ee16bd397c703565cbef54fbb4693b8fb1e48ba",
      x"0aa86c6ed7b2fe85574797d499761785b989133d37ec9122b5caed5b8e27e6d6",
      x"c9d3896fc3609043379b7935ce9aa001b9e5e1557af4b724549eba46d1aef50e",
      x"191f31d51470dfed5e3b1b48ad4d4cb29627e941e6de8aa54fb07ad1a9f73203",
      x"916586455b4c3997c5b14f19a1a503d677b47575201067704e8dd77e548adb9d",
      x"7e9d079d23883d42e1ec02f30979cd1c98784766a39d9a2a6622881fbc4fb823",
      x"223a729a8b06edd027f5389d3ee7ec8b38cb643e7ba6818a0defd1940ae4cf63",
      x"6afa7f1ab1057f3cfe24dec13e42819a5da5aa6e4d54ba83d07a264d36453e06",
      x"3e765274f263e917332d1f820ab851a4534122de8664798cfe557f32fcbc408a",
      x"cc4db1507d0c891d27cf6b8aaead20214b72590304dc97711492623754fd8404",
      x"793f66dcb807b4ac3d6004d4fcdfaebc45900f6489db135abb7633bc29081464",
      x"446f29eb26ec994fc3bf3902de0f3745fc25c0c1a8c3ff1577c548ce0f7da5f8",
      x"7628cbd456e7fd6dba9d72505a40b09343f751cd73739cd7485dae6f1e9e6850",
      x"43e3ebe55d6d5d801e139d74ae4ebb6a2adb2a1d4eebbc038f75bff1ea9c68f7",
      x"be3ed9e657669464e09e7770f590c0e6393dadf3ce995af69c5e5cf6312e50cd",
      x"87d19a990b058295272c704e83521e0f5ddfb4a56549e7ad9af077a8b9cc2b8e",
      x"5ad2e0389f4abb2fa3b2aeaa028651735025fc056ea20d6b62b0a499468571b3",
      x"5444197c7edaefc1e2f58747e310c52ef717151ae112c92870eef212f853355b",
      x"7b90f9193b7be4b36f467cbf6573e4f424968f9b077d626de479d9bae59f89a6",
      x"9bfb1e207f4bda788ea4e0fe8e376ce1a64d8643ec29789612b5fcc424fd33e4",
      x"5b61fc1d54b2a68d3245316df6f849c178238b927eac8aaae7278ff49d5de01b",
      x"0fbac216b7918a2b257817eaf77dc1545f527f14b77555497ccbbba2635f2f53",
      x"e7372a66a0a15439ccb15dd105e30fb64056b3fb9ec17b65b3dec28d80acce46",
      x"9071b6ca815097cd3f0e0382fc62dd72376200716f4439d93d19bfd1dcb73177",
      x"3897525795766f3999f43959bd43eb05b16e7c3b1777458a6cac62c43c40c8c3",
      x"495dad9482834a3f2b3dc37612f7eb53641e98701e0c50a6fb0717198de95aab",
      x"5268fb20282127d5f8d65f57de21fed4a7b3ebfa385d30d8b4623d304be7bc34",
      x"3ebc979a12c0cb867b1b7f298715b6eece8ef922fd9e0fae578fa17f076e22f6",
      x"9a5fd1c372c2b624a5a3468f8a2960367be0717bb7881b3f4eb0ef8955fbef2e",
      x"05d648f79dbf43bd29b73712b94b6588c78411071f508a269e53950d888c196a",
      x"75c965cbdbfbb2f2943c4aca1129d765b6cbd446c44cc27b306f015871f284ca",
      x"b332f27b15d34dc8a313f19c1599629a06f99f217668b372edc465e69e0109e9",
      x"e5a3d580d36df8ffb74174912e5996a4456159df4236e423d5b22c922f520087",
      x"55b3949082012376b2526b80f398a013946050276777f183900cb5fc1abc5f74",
      x"d40f1dccbdfa20f516c363d304cc0f448d6dc6b29cde5a5b91f038548033e3b9",
      x"1c6f1769473e0db4e6c502ca4c62c2948171ea618d3d7f35e7726ec254480aec",
      x"79290005477fb036e39c3f85051e2f611173df2d2217cc98fa7568851309d9b1",
      x"1bc4b1ba6b2ca788e73cc1fd2553b0bd7bcd9041e66d0828f4de0bd241bbe280",
      x"f587704c813e3891d0ed5af1276941a17fa735291c6bdc8ea689d81b265112f5",
      x"1eac4face46f05be4d81d618a37f3aff156d78d4ea0158ca0c27eade8276c638",
      x"12cfc6c438e2f69f551625aad8c92354f6defff546c0dc40bef8f977986e1630",
      x"67c9766a8d4d1dd5d5b32ec54bdf173f5e2e3c9e7f63eab058fb91ef74f8bece",
      x"e5d18c7c5f19e176675595338a638d3b1342329ac4e6846dd89ccbda6d4dcb5b",
      x"d0487f3bd86e0a6e4bc10d1b4af251a4a0bb7c21d08dc4b150ef7e5291011a60",
      x"3a81f7a95ca8417dc257a44b15c2579fcb545ce11a6434c97009aa9f209c3147",
      x"ddf5f080b2ee9fd5e38235beec76a24ecb79cd35aecc4846af07216050f7d248",
      x"83c0ae920705c0a121e5c010a3f08cea7eefcbbdf271f3fb99e0ddb1425850bc",
      x"e66607d02083f08978b8b97fd795bc50d2d38aa2430dc541335a79220816f247",
      x"e1bdc8c204d680956d94f556aa74746bea7fc4b775904f0e2208e913efa86041",
      x"9cad0914b69b98bf8eb0d48ef51fbaf298df05c34ef440e2e69272bd730e2459",
      x"98bbb191aa53b685fe4cac1a7bafd1ef3b3e1e03dcfc47c1bd62e4d4f3082c4e",
      x"a59f8f0f4f511ffbd2278d7a77220fb1d1a4722d5378b56e31cf2f7ba9be59ed",
      x"9cd190f5dc89748b2b63e829a311fa1ad00f8b33d29a077983018294854fb266",
      x"243cb5f7555a56ab678b74f3ef74e653227f1c04f82944fa7835fce9de4b5cf1",
      x"b843d40202e69153cba2765f579b1f4fe2a702c82bb2b529d1f49032669a59a2",
      x"eec053194f015de623dec91c3bdae831bc610cf3558414dc6141f8eb1cb70db0",
      x"a006c7c24e3f2808fc5a72e68fcfe4ec3909a8b711618b7932bfd40e4879abee",
      x"1bf5b6fb6b9bb2fe1df6a9657c637917ab5ea6abc5d48ff236e4f72ff8e13b9f",
      x"d125567ba1c1f3d208533eb047a9443a06805f2d46b80a5a0347092fe7812b43",
      x"0b8d3d114d2430660fa95a3a71c609a02f220e448631d919db8b0f2eb41b58bd",
      x"5c7461038d1acffa96d8b0db3ed998646e545eacd915fd99157c84ace62c968b",
      x"1717d09f8f84954d8d56f7b7daa9045164ce94a349eac15e9d12bd9ec5a75649",
      x"2ebfe0bb06718953784fdbaebb3eb027b1552b1a938b890f176656f71dbfd995",
      x"96ccbf86f446a149ddd78dd8b953afea74669e088b64feb562c2dc31bd0bb5cf",
      x"871e4dd31dc2ad1afb520794f176114fbe008615dd5a2bf01bd9f78456cb0824",
      x"f96a97a6b0b72bbf8d1f813a7be0003958f48f156931eef52eb52ed55cad80be",
      x"306afed323243fecf532aa958d8b974ec3b60fa344c851f497aec871f001cc99",
      x"31f5ec03be5deb1f46d1b417c4372362507e1608b9cc9995412a840bd97c4b35",
      x"4148afe02f112028a69fd305d820c37a221c0d3fcf3dc205039fd43f93017bcc",
      x"6ae8e268525d0de212a1671817ea04ffcf57dca53fd4ca4c8acc7fb81e424b87",
      x"6e4e30dbd1358ba1f8505ff2c4daca15565aadb5402ca4a7584bdc4055c81b22",
      x"dbd73b1258f47303eac6470120a589eab1d51efc8b162dd0a0d9df35436047be",
      x"297368a11649c444bf839af90d591ab802356b27127a3c786d86f79b3332fc27",
      x"5fa36199488f4034ff7a310e5cab8d58badbbe645500a39c760a8ca4535541c7",
      x"5cb016b16533cc869f721bf068678234f5b7b799608eb0fb301a575166042d46",
      x"f599409021004b538e82bececf01370a6cad301d4a54f1cd7a8bb677aa9a27e9",
      x"406b2633e2d042db284dbafa90ec574d127411b60336cb72ea0d4678b82985fb",
      x"7de70eae2492463939f8f52459bb71dbf51fc466455b1f8ea3038d6ccac4c2aa",
      x"29a0cfba39f9a894fa6e77e5487532f84ee7a2c4a4ab906982ab1b69da566d77",
      x"6a75ea66dffb2f08baa45d04db3e4f394b22e2cda9ca978fa1d5374c135bb0ae",
      x"d0f65e85f6c7bf34fe70e40f48552c2f4ae3e923df6b38679763508fe3afc0b3",
      x"b7d76045e203655410558fd39ed5b0861fa7b81da5b9f14067dc742ea7556fbc",
      x"9e50bab2477b8e0faa9a3d11ac08e690e62c814134599c47a342f65ba5470607",
      x"e654854578dd5b8e366ce6da7a7089d905523e08152703b1e216d2d0df3861f4",
      x"584388b7fcda7db36cfa2a50cec915ea0733eaad514e95fb571b1140febf0c85",
      x"07b618c24b7ec462684def3132db8d9688b0576b6ca30f46d59acc17fa58234a",
      x"74a1a25be5b8a1a369163f913d29de4256b2caf723cf55d9322c2f57a8f5008f",
      x"2da98be571ce34478a717e1ff2356934238a6615f050292cd2352a7ca08d430d",
      x"73a3ff76533067da99c3ea3699ef7d3855cbae2cf34be9bab5eb14f2d2ec59f7",
      x"da6fe2efb65dde3d5e112fc0f196cbee7b97b270a84078cb48bdef7a82a692f2",
      x"d1b984fdebc75bd98cb6595c04d23cff0e897f6279696a3ac1b7f0e4f2c5631d",
      x"7a8f25fc4e286ae72ff1d23056bb21d7a1fbed1aca25511cffb32fa6f3de8c4c",
      x"66fd92423c5a9be5e71509ae6ed7f5d3496c46fd3ca5caf596d6e32343a65542",
      x"f18156a3b0508a87bfeedcacddac02122e8b4038859294a6348966b0d4fcd60c",
      x"f95af991ee802d700c0a461b74d4cfadaacb63f59f874066777b35ce9cf6f441",
      x"8b892f911fcb086ab9f2b5659c3e88882e328c9d9bb27b96d6733897271b868c",
      x"74ead415d7ea9fe20c7bfd8e21ef1cb785c4fca82b5d164e8a1bbb8df68d1f87",
      x"8665790634948f64a95cac43c904227b808abd212bb41c7a2b99adb71c2e34eb",
      x"47ea07f67efd3623e99332c70e55486002abcede6e4fde2612f1b0c957443884",
      x"e25078ef9e6bbbd052951356547a045bee9d3b70e42a53084c990d4e0d3f5893",
      x"4166786f0054f20dd14bec27fd488f1e64d7c8e6b1ed0f46f553310db08701cc",
      x"e5d53fbb76fd4c5204536c17e78fb5f0bbdb6f396aa8ed7e7dd8e59d0a1ca91b",
      x"cf104fa25846532979d47a5c005f0c580cee475b16bfaf16958ca53a5c1333f4",
      x"9a2100aa1f82c2c08d0d6441fdcfe8bd421186a28441bf3d642900d677ab4b1d",
      x"0e39da9c7ac1ff351e79980c4ad20092594c91b66f15cfa9e03b308801c5f6e2",
      x"03031bb3333ee512ee391bad70dedaf979154535c5310232527f4d891e45e5af",
      x"ed4c76373d3467c7e2cab1a4e040835849344e850a6fa0cdebd478e898ad01ff",
      x"d4aab35a456b32fafc4ffc08c6a0d142871c53d4b2a4b92cb639bbd164647b0b",
      x"15d937db963f79232f785fa75308bc671c6d8f8eddecc256f7851e6db45dfbd8",
      x"f6fd8a27913925cf57f8e8523503b660cbcbeeeaa2c725eac1bcb9d4d44f3204",
      x"282cabfd5803cbbdf152713da9b33347e7ad9834e20ef1af7a33435756198459",
      x"6f93332ec3ab894537870e0f03356756377bcd5a683ae35bd8421ef0067b8d41",
      x"059014afd6b964e7ea2f63e5854d9b1886e84a1ab6231aafa00f991f37ac879c",
      x"483b8d2b89b6b6d0ec3769abe1602dd8fa77b28c216b28839564c07a0ad149c7",
      x"f32ef9153ea28b871c7f92b3e7bde60587e85dd753404d2cecb492aed2728a91",
      x"56bed236e77788ea7bb63d71296d2aec0fffe58bbf6047c05ef137d994bb6eba",
      x"d2a39cd70dfa7ff7b13fb065b8b4b216978070bb707c2de58ca3663e96ba7fab",
      x"27995c8f900e4b5a4d971b913c7e29c710f1b05e380472ebd3107071b46672f6",
      x"dc704ff341dacf1079d48b1392c2ed8415426dc73311c34eff42d21a0132b326",
      x"a07646ac5c3c17c03ebda9bf407f841c796d561d9cae00f3073f783d573f3627",
      x"221440e0b9944df2d20a66a3441094ef22e02c6fdc991554c6bac81a55a2118f",
      x"3e1ec0b9310cbd17522d3d34d2abf07ac8a56315611461345353c9b1bc98c63c",
      x"ef41c2ed81ef0a47605528d6fd29f5566816e8988df9fed85d157075330742b3",
      x"002d9b3f44cdfa3f520bbfe0023fef70417431c50634e61553001a057a6b437b",
      x"61c4d5b0ae96ef48bea47bae6d0ad5b140c3900828b44c4ca63b54fd3a2714ca",
      x"bf59fda1e5462f962d576f3bfb4d539ed4b075fcf5730110e84f79a8d9143f3d",
      x"06bd62897f212bd67dbab1b1eaec8f9e799cb24b6aadfb8b0e28697e4a085c72",
      x"7b6511ac65fef7f5d03b7c6d4517dd5893a616804548fd4c7a2bf0e978922711",
      x"fc855f84c22da97746efd547333626bd0a463471b385937fbe386d1839536413",
      x"972482bd42d1051e0a22480ef96df6ae598ec1471226ed890b044f52d12eafaf",
      x"6f17e205b449697206aed6586220e12a90a8ad8d98f524eb2e11f885b2b2c5a0",
      x"9f1b2aecb1faf828258c659569d2f570c6abbeab3a43e2e1b3173343fe3a17cb",
      x"4321366d750608820b66e71fdd00d4d102e269c1eabe4d116a8ffc76d090d4b1",
      x"0bc4b3843d0570776facf9c1b95cdf382d9ff51aa06be15354c9005fb76aba63",
      x"2bb2bd4d0f8cf356031da966a57daf88e0696d37db83adc6521f9c23c9ea84a3",
      x"106bb5a46ceace0af7e96d289048ccbc213731c8ae8a1cec81e8101e01b88de5",
      x"cdf1b95294f0e6dd34a83796c4f81bfe535d090537eb203022eb7c118d20b448",
      x"11a8fe9c329701aec08b21630a18925c65f87ed39e9c3af2c59ca2163d0a9287",
      x"2336fff5881a3308a304884b0f981df74330634e3fb2d7fcebe3fdb974a973f5",
      x"49b1f1cfd43a547f58793a7a8c6dd22f1c6a907de4c0a2dff25d55cde3878ba7",
      x"879f8cbb25751713be85693b49c78690bb010466734d8808aac06a25884bfd9a",
      x"67f61673d2bbbc734d53b28da6982e4a3366191a178b3631e079c78662ed4fac",
      x"002e79a42691defe88000c75b6f63d45af0c0c218551e96fb87d5b713ca377ad",
      x"39e64a1599bfb60268313e4d5efa3dacec910b4e2fb77c2eb852687b2aa5cf9c",
      x"9cff86d88a75f800e5f696ffc827047fec2d46d4061de25eebdfc3c7adcef65c"
    )
  );


end lowmc_pkg;
