library ieee;
use ieee.std_logic_1164.all;

library work;

package lowmc_pkg is
  constant N : integer := 128;
  constant K : integer := 128;
  constant M : integer := 25;
  constant R : integer := 11;
  constant S : integer := 75;

  type T_NK_MATRIX is array(0 to N - 1) of std_logic_vector(K - 1 downto 0);
  type T_NN_MATRIX is array(0 to N - 1) of std_logic_vector(N - 1 downto 0);
  type T_SK_MATRIX is array(0 to S - 1) of std_logic_vector(K - 1 downto 0);
  type T_SN_MATRIX is array(0 to S - 1) of std_logic_vector(N - 1 downto 0);
  type T_NSS_MATRIX is array(0 to (N - S) - 1) of std_logic_vector(S - 1 downto 0);
  type T_RS_MATRIX is array(0 to R - 1) of std_logic_vector(S - 1 downto 0);

  type T_KMATRIX is array (0 to R - 1) of T_SK_MATRIX;
  type T_ZMATRIX is array (0 to R - 2) of T_SN_MATRIX;
  type T_RMATRIX is array (0 to R - 2) of T_NSS_MATRIX;

  constant K0 : T_NK_MATRIX := (
      x"ba19e4d0e3ecedbbaf6de2130db3fab6",
      x"d01f5f13b96e762cad00d790bd7ec09b",
      x"66f907cded493c06b637f81d50777b16",
      x"aae722b6883a480acfbc1f24785efb83",
      x"a24778030fe971017beee0d6ef1be8e9",
      x"d7613bdc8b0db3ae6babec0353cfa2cd",
      x"74b11c7c21d673646ef3447bc1548d35",
      x"2c523cdd60792a89ecf4ce25a6afc827",
      x"595a780f3ec62d3c31c85941aa703c97",
      x"575cfc912f9b23559211e8a6ac31c63a",
      x"fba479bd329f29fea8b875074b3f3bcb",
      x"98a0116e68f53d5ed3688070212b96b6",
      x"756d45155883793e4ada492524474849",
      x"af5071ab862dd445cde52290c77d31fe",
      x"26c36753a6a569521c0ef76eea16eede",
      x"9a83a95b317bd6a5e2fc2efd4790cb29",
      x"88fa21ff56c4ad3c6f22ecccf290a4ce",
      x"60b108a897b009fa1547c851273e3c39",
      x"f7e3b742d6b51239923bcc725b6ef64a",
      x"c6047a174d25cd5ca922dfaadaf3a3b1",
      x"ba904c992f6342a55b7f58996ba09a28",
      x"50837e1134dd246331028ebf5b543fae",
      x"6eff54a066f08e9c38b568c389446549",
      x"9b26aa662598fec46f9fcab0dcf2de8c",
      x"e322b0c557e4c4eb2f36e76d06c8758e",
      x"76a7a3d92c5527ff4bdbb39ee07d0043",
      x"6822a366b640284056889c1af1ebe56e",
      x"3c55c3e8bb148980fca9fa272064653d",
      x"acc88848700190126e4fc4ff96cdeae7",
      x"709e01e10ecb01cb8a1abf792adfaf2a",
      x"0bb94d002d8335e44441310499af1a39",
      x"9363105b59809e25692fe392266b1df0",
      x"2412d12d9866b3628afc28dd30eb4eae",
      x"5313abebc094f0a143dbd3dc6cdae341",
      x"1e4e443e404e6707e6a7630171f54507",
      x"975a09d7711fd32cc6e9dd93765601a5",
      x"38a30b7b059f9ecc418745d61198afee",
      x"8814a89f6c5437a7e66ff05f69ababbb",
      x"f2cab6de907409f4c4f45dcb6da933f0",
      x"95a2ef55d78091207c824babaa74e906",
      x"0bc4f487cc3436b8982c9785d2e75d5d",
      x"74da8347f644563facc56f7b1455e8de",
      x"f6dbf281c1ce8ddc71b8a2ca331135b0",
      x"30634eb239fe2efa72f46249aa3fb300",
      x"0214d09dbf071655c607426e34f72c39",
      x"abbb61b5be7262e4e2e4b14dc3c2d08c",
      x"e6e55a047828cc8b864d7a6b602ed26c",
      x"7264bcd6d5c82b78131034167f55f40e",
      x"36398b447d98b72bce83f6a4de5d2840",
      x"7e99a3ff909432e871ee4b4594cdc032",
      x"989723d685f60108b088e9b8962fd824",
      x"979e6edd870af0567efa99d5fa722a2d",
      x"da03d220104e0ca9b21093f28ae0e65f",
      x"c255b3c63df7e7b24192582697f3f922",
      x"ba6d625959c5d71e24b8440a26003c0a",
      x"e419f3f2cd4d454457d177807d6eae88",
      x"9c7ff8c5a55b195eebf51d162d5fa682",
      x"bdb80d3189ce779fcf3d7588009c48ae",
      x"b68356d4f6b2635b766dbb99ef5fb724",
      x"284fef4881e65d8a8658c04cdd78f129",
      x"71164bd236d0a6638595cc41f99967b9",
      x"396a2f6246b3662d486ed0c5de0b8e7a",
      x"fdb3b984a81fb97ba943af45a27e52fd",
      x"62846cf34cbf677a74bf1288cad67d99",
      x"a65bcf3d97282eaf19228a007fd23a41",
      x"767379feabff651e9526e8dc04da8cad",
      x"504a980cf0c7a91d7df6513101684d83",
      x"d24dfe828f15467fcbc440deab638e5c",
      x"11ff4f98c5a638810d95fb4d3fa79a59",
      x"fb81076a6c99d87ca145d9d43f3f99e2",
      x"4261f8d834f3010451b4d470902702ed",
      x"3bc65904d54f18e846c76d32ca0c3f9a",
      x"4c749a851ed8a794d8742edfbeb6b75f",
      x"32aa73b5607c58180bea37ed2b16def0",
      x"8f278e34e2a392906c51fc68045582ac",
      x"c82fded0e5cea98052ba63afac3f7870",
      x"e833360e2c5c627e7ce509b962782ba7",
      x"b670dd86a0414be4fa2c57cd2ba88589",
      x"7c56a83fe943c97a7d6d092203812301",
      x"8e3a1b85b05114c7dfe4c7e6ba0846e6",
      x"1815333b6b341a0631d53fa11966f842",
      x"2888f850f91315d83fb762b5c6314915",
      x"035f429132aa6d8ddd8f22eeca228a3d",
      x"83f9ffd7a0af3fa78e00769b65dade57",
      x"390281b53921d175d519ce91003e6037",
      x"2d8559219616fe4bf567048e7ad04b11",
      x"e22afb560316d4000fc50744c54731d8",
      x"92b61d1607ccd28d5a752598a0d15bf6",
      x"e16054452053d05d3ba20b181f47c519",
      x"03cef89085b4ef711ba36dea0630285b",
      x"8376a952fa46afff0eeb600170355cf9",
      x"b7b71df107a9c2937a7be1d03047bf0b",
      x"20f4cbb58ebba98022c3e3dc47993997",
      x"055a2cf1003360fce77a60f6092b09ba",
      x"8bd192d49a9fde7a76b27c1cf22e7e6c",
      x"5adb106693828c33134f671132f6579f",
      x"a2853c664e3153307e899da03c1b8ae4",
      x"3bb49336c2fb2c6e6dedc30083e52c00",
      x"ee4ea6975a9eaa318e2fae513306ca91",
      x"47f236715c5dbe72a5ab6129f79cccfa",
      x"d6eed5d90f247ec1a7ef7c0d704cb6d0",
      x"6f1bc7447ec7b18562f1d7e624accfba",
      x"59acdc0fc574e96720f808e781057ffa",
      x"83089229fa37c8573d9ba780564fe5af",
      x"eba55f55ea11e152a7870d34abab319a",
      x"cecb60cb456fe77d0323ffe9b05b67f4",
      x"d7dfaf3a880cbde6cddf331c6e0f7d09",
      x"b799a351be30f819f786003395f8c6e5",
      x"10459758c11ae4849d619bede075362f",
      x"e57868a81ca45d60d9abf142dfe01b2e",
      x"c925637529736b1f520607ed73860f9d",
      x"f6db108ea53663362b42faed50176c0e",
      x"9442fde0a1d42614a55ad2a6dd2362c2",
      x"2a9940c79ffe32a6aa4c6d60a9fa8db8",
      x"a797dc31d0657de1fad0e9bed3db7ae0",
      x"b5c51493011ffa691640e20ea18dcf02",
      x"40aa4ccd7ff48582901b3053a356ee13",
      x"93726b123cf09dadb1c07b2b2956b138",
      x"2317d2baaacd086a72d77cb1f81f3278",
      x"99aeb29605ca8b084607a428c08ce657",
      x"14f72a5c66c81e7b07fa92c8f451a92e",
      x"b4983ddf65ac129256bba0118a7e8dcd",
      x"38aa769e34b2aa11381f037048131cc3",
      x"d4e102b60495a28d16515998df284028",
      x"be44f5f9b81879d5c333571e7988b510",
      x"1011a19f789685084f7f1459426c338f",
      x"5d0a069fae5127a15e58b761f83419fa",
      x"289fe961dee3050429a3782c031c443a"
  );

  constant KMATRIX : T_KMATRIX := (
    (
      x"b4809fb0d897847f7b6b51181b914190",
      x"057b87b942a1e798949435768b05e66c",
      x"43544fe920fc6978e074f19d5af2fe3b",
      x"ce78553746f1498adf8519b35fdce812",
      x"51d7403a31bd24cc643908212092b04a",
      x"18580c3fdbd709e6a3c405aafc11fc1e",
      x"b9baed10939a3a6a84d7a95434a97cac",
      x"5bf05946f4b1a235e7a647c6dd74ab2e",
      x"28e643c39576db2a219a69060bb2cd6c",
      x"ccbaf1a931680ec0c884c486674de8af",
      x"de361f5b9c5c85b3f3f070762d897f9a",
      x"2e837a3ecda13f3efcd791db3ce29d70",
      x"f37960eb5fe16040889ec67e8c2a7345",
      x"af9727cadf4dfb8c4a34d276ce4620aa",
      x"0d2787a7ae5b5d59c044b047c200811b",
      x"b581740379e9a39174636848b937fb79",
      x"b0840db3661c0e0932f81e252cd1311e",
      x"880700859b78505fb88f8ca56ac918c1",
      x"3699d3644fb47dc0291516b4b828a16b",
      x"ad3ee505e37a16042056cbb2d1e81242",
      x"9a0e1609a7c5fc2693e133b7316b9c7d",
      x"a9f918709be10ea73371392c612162b3",
      x"af458cdcfe83bae63a2e731a2018c758",
      x"dd81bca382e802d609cb7762eb1df1c4",
      x"e1d6cb27b5992c073210909176ea30a0",
      x"453c09ea8c07ec400ebe346605540908",
      x"714a9f46972480aad9f8306bdc30721d",
      x"7fab8309a382b012cd5c7eab2bc57f87",
      x"83ef6e09649b90b70384fa7dbe03ac3a",
      x"b703e1996920d0c306ae8265f45079e1",
      x"596e55c37b6e1fc95b4e7fd6ee1a8958",
      x"a6ce90f7f4ea5b754d82ec0f1cb4bb84",
      x"226f12809bfc27098da7773f6bf89458",
      x"a69223a469f8e3b29edb443712d44959",
      x"62acd26084714aab707ecdce76db7afa",
      x"31e571bf5ff1b7f19c361d46609370cf",
      x"0fbb2a1aea6f81890b1ddaa4a6b88ae3",
      x"ccb484eeaf0409146af9fea7fd1edde3",
      x"047067aee34ecfebff8c3673ec414b36",
      x"59b13de43673ae568b1a432cd2e31e12",
      x"cf793228dbc86c334065d52f9e99168e",
      x"1dc791f89342d0d19a84202910e64adb",
      x"4238d1c3d23dd037e6876f9d106b745a",
      x"1a8d8cbbb8674f3c1df8565f0c4fbabb",
      x"ac75b855c09c03addcdb4e9a433f2084",
      x"7de3e55f3c0bd15997162932a44716bb",
      x"139988a2684b7e12e621529648cee4c5",
      x"eb39df8d4ba9fef51c70d0aaa541b15c",
      x"8d484276278653a082b61c3779bb31ba",
      x"3fa975dae7c25f49434749483442b796",
      x"9d104b69fdd0eefde9a671bde1fdf0e6",
      x"de93e94a95995e6704f4a4c333e3a3ec",
      x"9f3cf2e5156b3538b4e564249441787d",
      x"463ce0c44d0e509892e106e7af7fbab5",
      x"29d04b1f08ae22abcead64b39d284d62",
      x"277764435ca5028ecfc843cf3fe96c11",
      x"8babfd37efbf63796ca0a72fbf9d0334",
      x"cf6901ea7d310b978f101d3b3cb1f172",
      x"943133176c392e2dcfb808de22c86ac2",
      x"1002279c17ea5e67cf2f4181598e08d2",
      x"18531a33dde27bcb4e10b98663d08b3f",
      x"74f002a75e46df89f34191baeed868c3",
      x"96a7f7efe024be42fbc59d61fd902b93",
      x"5035c912b88bda3c80a688aee7fd7658",
      x"928a85846d6a519b400bdec7251e8ff5",
      x"e1c50906337f18b687a467d9e9a0f071",
      x"eb4a1c5cdcd1331cd5e88b6187cd33dc",
      x"f6edaf4c044bf619ed07b0749f370c4d",
      x"b9bc8ca1c58b8ccc85af40701eed51d3",
      x"c906a2f40de7a949e1c00ece238072b4",
      x"df32e19f59869773c7e983c3b8dcf96a",
      x"3f759450eae0da487c9717c153f22655",
      x"f3c85e3c20ad6c97878d43d6302164ed",
      x"857ad54fce64cf30b8feb67e9e56882f",
      x"094d17aca923c8d6b9110c4138fb6276"
    ),
    (
      x"2488f659513e25fc6408b0e0ad5cdf9f",
      x"ab85a3ed46ea5d78f99a4c417a2fd351",
      x"bf397e0e1d66e6f499d46640859449f1",
      x"fa15033430cc7c0d271ce09de1f2535d",
      x"ea474dc408008db9f6460f5b9d5d2bfc",
      x"1859db0390d9bcaeb162e639b3bff380",
      x"7288e2a16c8a09da0c6f9e2787293052",
      x"d5f05227efcae364a2ac5f513fc62602",
      x"6cb2dfb90f2c58ddff61e36877e7a352",
      x"559b04ff09009dcf67662519f38b2171",
      x"f4c08518ecafe3260d959047356e96e4",
      x"58faf86bfa13b8a40ee2974e2bfcc8e9",
      x"7abfce5f770a31e702646f3b090e9846",
      x"a648b4f299ce7197f3a68570fb6ab6d9",
      x"be76bc097251c4d291f34e6f68cf77e2",
      x"a543d5c55c8db4c633aaef6102f3fde9",
      x"938108106834a3bf4723a7829b9beb24",
      x"3919ce7daf2c6348342cb37778617e01",
      x"907d1a3fb9c739fab2ceb3d0cfaf671d",
      x"0490e4f7e51934a704b8c9a7624749d8",
      x"175c93f044b4841ab72636cc4c9ad0b0",
      x"8bf5e1b41601f7ebeab8af933f079de0",
      x"65fc87c640771fe9cd320b883093a00c",
      x"d325d910e5c6175325f15af726fd5c60",
      x"3282978ebae1ba4927c1232f9d125792",
      x"b154e966e00c964161a81f53a328953f",
      x"f295c2d91e9099bf969862a16e242393",
      x"0c908432f8ab39964f0dd51debb89960",
      x"fc4769036f370600c7dc175d7049ea8d",
      x"ebcf8e865a22122a2b26d333b02ae45f",
      x"f29796c493eac9918ea469117e380d21",
      x"1868cd7f66d168e43446828a2df29857",
      x"6a54e87d0f4c3ebe692d28dc551c3fbf",
      x"132bbe7fc3c681e5680cb93c3c27a75e",
      x"e09b77f2378fe7597fde7eeaba510ea4",
      x"97b5ab2f60fdb72d2327af72a4905ddd",
      x"b27d2502596466b326fc4a7fd662832e",
      x"dbc6507331722aa1acaa6d6c42098f9d",
      x"09f420711bd52fce5ecd7b6e41b740b0",
      x"bdd7cab939de841a48c6e315b79890d1",
      x"df296824d704f0055b5b34beca7a0996",
      x"5cbe3bc6be63891a298c6667dd907dc7",
      x"0d28ee9374bbaffe60df58d02c611440",
      x"84b808f79eed45afa03a1ace733684a7",
      x"e01d05fed2cece58ba752624723525eb",
      x"31063c6e195e3dea24ff72ad60570992",
      x"e3311360d85e7c8e5370d4bfbabd817f",
      x"9e0e36fd54149674b43fe3597e00ba21",
      x"02c4233df5399f8c59906fb400f92878",
      x"6d568bbd5b5ddfefeadf852796480a86",
      x"e9f1dc2ee69222cc5fa4ebd0fa2ddc9e",
      x"1124a7ba5f9020d8c54e3158b5332c49",
      x"f97df25b0c178868b874418c229cd9f8",
      x"17447003c513b7b5cefdf9ce77e85063",
      x"d15c844548366c921c5134acddded8a8",
      x"cc97c1295a61d3fa83c5a0ab0f5f3e47",
      x"b0b17dfd1815f75e7d577d305f2bcddc",
      x"c9499a5bb25d704a2d13c922b3cb917e",
      x"e39b8537fd0b67f89a5aff9025d37fd5",
      x"ffca7c11362e5afbf8bb46e30f4ba5d6",
      x"d93b391399fe994f0fd561d3d7845391",
      x"f4d1937403d768ad45eb177d4a1b881e",
      x"1a3f42981078355b2a71b373c1731610",
      x"cc4b07c2f9a598759ad2693fbc951d76",
      x"289fc974dbf2670d2c5a72ea274fd305",
      x"60f767ddde9173afc7a1454f15c6fdaa",
      x"5b104790657dce73c429b08c02f76dc4",
      x"2115c0f81bcfaf691fcab05a7b190f83",
      x"eb8df8a494d8724ed52e5f5e42303ed8",
      x"8d96fce936767ee54fbeda9665e55183",
      x"6cae3de47d1b2dc1e0f89cf6961b6abf",
      x"e914479b433a3e3b7c4b41f091213799",
      x"1ca3bb55a9dee16b79fd8d2660d03bd4",
      x"1f4c776fb5aa9f6baaf765fd00a832d7",
      x"e15f76aac106442f49a9bd58739a2efa"
    ),
    (
      x"d4cbeb645be809c3d4b275dcf10b38d8",
      x"5cd7b1bae96c64917e05072412698c81",
      x"de0f550cfe6414fefc36c0dc2ac15cc2",
      x"e5f5cde7d375213bd77c68429ac78d70",
      x"0ec5d0496d24eeee64c997667176a336",
      x"bd4f2576dfd7fa7e71cfc7aa7773fafb",
      x"5e418aff7e9a7526fb4fe0ada8e682f6",
      x"f783c7152c6acd4e96d216002bc41618",
      x"2bbb1952ca19545859b6c5da658cbd18",
      x"b5963fc02beae9a9a3af22da3d1f8efa",
      x"be3e4d85f7a6a331336b9f486db11e5c",
      x"87c4b1e60967c13139aec4e26a0123dd",
      x"50d010bae4ac215e9d564cb255aed775",
      x"b820f4e57f0fed37ec047973b59cb3a4",
      x"2374b2fa454ccb5977dc9df8a7bedb48",
      x"cb7e5b7a19989694a0bd5cbfcdf329ac",
      x"4edada96c06484bbd2eef48525ba6949",
      x"b8d71580959a7afeec5f89567e252826",
      x"703d4e1dc4ffcfe26d3d49114f560741",
      x"711c260cfb9b8bdff53ee9eec545166e",
      x"cf28171c46a6295efbf17f694f90ecc0",
      x"75b407813aa3660d0a6ca64a8f24afd3",
      x"c84a1a22c70ce1be394e7907fdb5ccc1",
      x"c276fbafac12247e32aed3536318bee5",
      x"6b2b50a61184f374d6d0f8794532e665",
      x"70b7c3492d79a7bf178835650cda4e4b",
      x"63f54f6c98711e6ab2878a9a30b36d4e",
      x"926af23e57234add35327d5592c6017b",
      x"b663432e8937eb80e6efc66a252abef9",
      x"ef5c2fee0e05fac398f00c6ac4db7d99",
      x"a3a0fb21fbbbe903fe0a7e0e9329a841",
      x"d53e59b9cd1e7dec51427ccddba3012d",
      x"83e5524c89dfc85102362471920d4b54",
      x"db2a5440e26044481c18838698bc607c",
      x"c203fd718d7a280f4d3bab8f3a714d21",
      x"2258713f986e25bc0dcb6de26b736119",
      x"7e7e669e39f64b63b8de64c1b08b785a",
      x"eaf8388b64cbf62aa9aff01b5a2fcc26",
      x"7737d1b1beb245c7c8066ddceed64d84",
      x"e02c8f838bafab968e2cd64c9064dd5a",
      x"62e9f6142f2b68db1c0cd1f6b71baf0c",
      x"9dc930a490150f7ee830f333d0fe56d4",
      x"9b6443cdc8fe6749aadcd05ecde6dbda",
      x"756df712bd5bc19b97f1c102ce4165e0",
      x"5e51c2dfa0c945882cd77308348b5b41",
      x"7c0123ef7504473cafd2e48be3acfaa8",
      x"88459cf49ef26c463837f0759af4ac7f",
      x"22a81ce70b8c682805928d91d40783da",
      x"8a772dc7e1a42b4756eba3b065f420c7",
      x"8d605ff766da802a503210f5c137e537",
      x"08d1469a823540529255e8ead2a7e974",
      x"37bc434e5b47e5388cdcaa9a0ab959c6",
      x"915817e967672e08594e40e9e9c761b2",
      x"d345ed218a2835850c70c0450f7e30c7",
      x"be4086da86fbc27bc1c1ffa1d959f1c8",
      x"c733fbce6c06ba891e05a9153caf20cf",
      x"6022dd96a572c282c3b175796691df54",
      x"7a15a375e6a611b3a4d6789e1b21020b",
      x"14257c84479e91c72cbd789b3ad8ff08",
      x"6ce5dd6cc12589e22006cf6963545956",
      x"d87d0b67bc1f6bcc56b21b79fe180d16",
      x"757052206b91ee4f711b33fd7c2b1a65",
      x"c153d700e807a58aead1164bb8e0e9e1",
      x"24ac62d3a058e8667ee57832ed469a8b",
      x"1cf1aa39f52ab0b6de7b9f3989cacce4",
      x"6ea9ca0ce9fe0587a1db17014249dd33",
      x"1b7479ec4fa1dde3561e6dea0bf5daae",
      x"e7d68017b1a38275c6b59ef6c9120f6d",
      x"a22bad605494c654548ad4a79c09489b",
      x"9d38d8e97b942103b4547fa02ecb3d0e",
      x"d6c6bcb554a3df46e8d3493a4bd6afab",
      x"ea5dab332672c2f3ebfa82c102d78154",
      x"61361e488650b77815a2f6e6c4b12afe",
      x"b4b1cae4f3e677ee14d3d5ec89669283",
      x"47ac4130fa44274fda9f708e31260a03"
    ),
    (
      x"35c35e2e372006b79920088d5d03c03b",
      x"35e6794d384328315dac3fd14ddd2904",
      x"b1d13108cd6e42ad105be67fb371cbb3",
      x"00b490aab382b20d3b1886cefcccd662",
      x"3d16011555c49f1631b1d6fad488228c",
      x"5814359eec8cef665d82078800b148a0",
      x"d009ecbd866a0c731bcbbe4841a87814",
      x"99a94022f258b00ef56d6c0a449daf4b",
      x"25a168e9fcda5eb9f6ee4aad0650c1e1",
      x"f93fb1a64526d6c4a649b86367203cbe",
      x"5566c01b2effc77291b383a0142b4d88",
      x"0733ea039977bea9116a527205118be1",
      x"d3995dadf7bb7bc1bb92b8a5ceaa9e72",
      x"9114b4caae6257aef6f897800619dcfd",
      x"f48d7ad027e11ca10cfded7d67e61b41",
      x"abd036dd81df3802dd97514f475b3406",
      x"a98dd9f098fa7eaae4c346be85acfd4b",
      x"2805f05fad368e7bf46d37df0b083ab5",
      x"2a2f112e6ae9c1ec9ec212d06a875a2b",
      x"dbf6608e69b074161c51f4c3eb59e593",
      x"911173b25a6c82730f740b09afffa867",
      x"0269c2c414a2ff6e841bc9410749ff15",
      x"b8a2d89c68132a2fb4e1ccdc2b01eff5",
      x"f2a2d1c1023876a08148013e8322247b",
      x"1d84f3e4cede2d14dd8c4bdf14b60e4c",
      x"93a37e330c99abb92c59fd2ea624b6d4",
      x"bfd9b4bdeec70d188007fb76ccbaa260",
      x"6f1ef75cad7b1bc25f6c15bea5514311",
      x"410b8a45ca51e93acccdf254b5c87299",
      x"532156ee0f8afb7b231bc9f0aae02513",
      x"b8c79fe7f2cbe9c2a7dfb08b492a9622",
      x"3e6a4b4229717b8447dcdc798b3fc26e",
      x"ef53c41a02691b28205429cb26d5edae",
      x"0e2eacb75697fbc770c7f0284eb2ced7",
      x"7efdada7e827b40ea8d6259388a70cc4",
      x"68947dfa7f99236ca95a4114c09d4483",
      x"57d74cbc1c47397ecca73fa539d1b068",
      x"9cb1b9124356d2c46fe17b39f8810d91",
      x"83c230a1fd1bb4194455cceef5b9ea4b",
      x"db11371c9e07be3c5718612410f4398b",
      x"b7ddf3bd9390eaad21787ad3a684eacd",
      x"6cdf27b42413b247f9a3c53ed387935f",
      x"2ab6023a3b67328f24b448ba23a7304f",
      x"beeafdec466cf65e8b294a8651a2145e",
      x"d06add4d8050a80cc4fb44d1495b4f14",
      x"29ee5ae7c97d2267f0ca9deb38cd73b2",
      x"189e5936da1a8296c169c7b62a57acf2",
      x"8bb3332a3338269f4da8bdfd7274c9d4",
      x"46ad9ba7f82c6c7522445cc585857d7e",
      x"c1df06525d44706807cc08413da68528",
      x"aada45fdd823548feff179fd58c59ab7",
      x"5510416e3857c33a624c65282a859c58",
      x"a5365cc0035a6b32de4c59f2a0f53680",
      x"b0a4333e5ae4687976d78221104c6f77",
      x"cadfe787604104a84a60ec4b31234e4a",
      x"fa20620b41e5b77c40a0407c8e25d6b8",
      x"9681993d130b62211629246250549bb9",
      x"5381eae80ff5b699fd345fc80e3c85bb",
      x"0b7c68f8e8de98969a6d9a8a873b435f",
      x"1324e01548c4a6e9ea5237ed36f21039",
      x"077c6e35238e0504810a434297b54fd4",
      x"ff59b4ae5209ea000a28d07b8b9380db",
      x"7bbae16a479ec07ba0e4b1abbcea5595",
      x"ea43f3cc6fdff0a79af0769a01643873",
      x"392e5ce9c81c8906a8f48cc3aee4be6b",
      x"43e29a645e0e6cabe0ddfec04ae6401f",
      x"ef3ac8a20e5d5fd9b99cd668aea46117",
      x"698dbed3895d629d94024a5489e038b1",
      x"ee9b8d636dd9a2c70faf48b34c7515ab",
      x"d2d0f77495a732cd9dc6c87eb8ec971d",
      x"e9c9e610db96283ed0bf0c8d06e14a86",
      x"4a2baa0af95e53dfcd5d9c2c9e5debdc",
      x"9c6966b1b3cb87c2eb009a34c69eb37f",
      x"551a19bd1037ecf72130ce973d981749",
      x"6e7311edc91138b643c7f778e2374e5b"
    ),
    (
      x"b854e0d45b863e51d2005d5f9e43f518",
      x"d968a414d21a6d7d45b34b2620fc7a8c",
      x"2b83b2499318f06e60bb18cb3873a4dc",
      x"42936416f27e1e8f8a362591c7256e89",
      x"f7fbedf3385ff49284da44ecb6b5d6dd",
      x"56e7e85e5b075280afd6da84ab42a5ed",
      x"6155e4d1b0bcd652c89dc42d4728fb31",
      x"7f91adddb76176125203aec5bd500481",
      x"41ba8de2a6ac955ee2a550fa09c35441",
      x"8c59adfeb5ee1b5774e4daef07b3752b",
      x"8bd40f59fa395ed406e653f9b6aaf272",
      x"8f78ecb7bd7099bc23a9831ec9f1cbbb",
      x"f7ac52e81b63fa5add2f8cadd07e64f3",
      x"cedcb226c9a8ffeb8f7a7dc4cf3262c4",
      x"fc658d0268a17b3acc82a5d09c28e435",
      x"a481085dd8a70a6cb2dd9ee5547017e2",
      x"acf13a35522d987e0cdb74293f400248",
      x"b7db0838285e4d505bc45d3a8c7451b2",
      x"0e097254747fc89468e1b9b79734cb0b",
      x"55a977f7189d02cd2aef7712d7697250",
      x"f3c815b4704cb4f4352107467fa8cb56",
      x"c44f883aa692272003a810cfd1277259",
      x"435454826ae2c893b425ebe43c79f746",
      x"943b2d64183625079475fa8261579a46",
      x"87dba33a8919ac293efe29da0587684b",
      x"6d2cc19a92d983dfff3ce65beed5630b",
      x"95b7a2327110db8b641ec433021dbd35",
      x"1e2298d316421c3d03b6f87b523eac9e",
      x"7e80d75dc84f942542371cfacbe40854",
      x"3cfc694110c46f25e9dc5ccb3de513ff",
      x"e103caf90c5ecfdc09ea57086ca38afa",
      x"d980200218dfd8f66426a1c7e7856352",
      x"5e812adf4b7a0835396ffb1223fb2989",
      x"dce64755623d55aadae0260cf37a04c2",
      x"98043bfae1934c2f72edbb1cb86750a8",
      x"23610a2705136a071cddfe6d09f81471",
      x"7632de272d5786fd2bdc81b2b5508afb",
      x"d2d233d4aae56b1bdd12b76294acbf19",
      x"a3334db6b70ba62e07a39a4e4abb8edd",
      x"6dfd3c1635159e1528162abe4d83a49c",
      x"cf8cf6d994affca62ce6f8053d6cb2c8",
      x"6a7d2e16590e009e3bde0a2b198113e1",
      x"935aeb86e95d2531ae7120c5ec57cde8",
      x"afdf935ac3622301364bb36935d4889a",
      x"9ad72a1bdbf1e7a108cdc861c7d31361",
      x"bce3c91bba9d989ffe5ae3772e44c0ce",
      x"a0900cf5ecf1da46b9c35860c76c9f78",
      x"3a963abefa4765b62bec29685399dba1",
      x"a3fd54985516a22d2d2512c088e07880",
      x"b7aec4b95108adfec0d71cd02116b1b5",
      x"671bb5416e071fe5b29fdcd6d420a79b",
      x"ab7f39318b700d9bb58dad6064c0a336",
      x"81de8c3d4c1c94964c44644056bbf8fa",
      x"71d48b08c5fa5dc5033c3a0bfa1ffa4a",
      x"12851733ef88bc99cf4b5dbea1ab27b1",
      x"b5616537f7a41d53168a941649726873",
      x"2041cb4b3c49a8049b20c91301deff78",
      x"6dea467bba8533760d56901284f4fdfc",
      x"708888fa1ed82c8ca843f0025edf2214",
      x"0577f957a533d7c8ad89c92661259ff8",
      x"71a568f93635ec81ed53831b629f3cde",
      x"8371a6e58bbaa11c5a295592436bb222",
      x"fe80b12de522b05d0db7e5b075ddf2cf",
      x"aee03a766874d6570f5c117a5a143f7e",
      x"009e74e3774866c17eebca4c4d93430e",
      x"ea485d3e5768ee9e1c7c05c7b91fe9c3",
      x"f1157026d1f31391b883c2ad6b31b5fa",
      x"da2fa846ca8774c62474722641759461",
      x"21d33f2629d3ef05db5110d23ac18ced",
      x"af6d88b78661d06d0b24ae1310f3f0b4",
      x"0c1a1e0efaed596306eea11fa03f6b45",
      x"2f65e8b343f84b4127d09705097b207d",
      x"260f9bf17cf32514ea700de53b171ee2",
      x"c7b76ef697b57de80648f4798eb54f67",
      x"18365db2700a378aa9dba34f78751920"
    ),
    (
      x"129b62f4a28e39ab77d328db4d77d6a3",
      x"9e8c72bc17d496b15f030e41063d85da",
      x"9993c36e931f09c075652395d4db6c81",
      x"283780f1b6e9a6596be7833051426260",
      x"90ab4d304363cbfb83c3dd4296c3673f",
      x"c7095d2717816a17f6f12581b048ddaa",
      x"35ad720c9e7ebae733028e0c9f7ca74e",
      x"dc3f731fd2ab45308ae1cdff62da7089",
      x"e7a4464fbcd1a82f53ae8a6f8a888fa4",
      x"163f3c8e03b6f9a78902c7b14dceb04a",
      x"e265e35a7ce907c4ca0f1cb2f879a402",
      x"1b331b2d9e53a029fb8644b5b6b829f4",
      x"998a5008d05183fb96bf9cdce153aaae",
      x"3f4861896ff3b02806ddda8ff442a327",
      x"3bd4c0c65058feefad95bb06d99258ee",
      x"dca2fcdea67eb6a72881a0ac5c635be2",
      x"46f85a5bb721c6a6404b073cec8720e9",
      x"90350df1bbc70a64033913c7f8afc5fb",
      x"8a98dacf783d9fe2f2d9142e23af8b91",
      x"0c253ea435012bb9c25d33d445853ee9",
      x"a349bfe4d2a423554f8b08ddb8984b4c",
      x"bb889ed7a42402dca5ffd4d8ac8bb5aa",
      x"e739c3daf47f30d8fd23284cdac08278",
      x"64dba128fc8728be62eb02e1b0b1fdee",
      x"8f4c766fe49146d2e17e98f46d4d503e",
      x"3c9ad87a1bd970c10ba38822f72cea7a",
      x"bcde6a27078565d6312876cb9a749c67",
      x"f2073219e9659306a43bbc0ff07b2784",
      x"65a7f1aa5b447c509c6dd868fa67b331",
      x"15e18ce2fdc17d12ff2f68b631bb1017",
      x"23ed8a8b7b7edac80d8904938996debe",
      x"0ea2f59b5e7a8eecd5221b77d573344e",
      x"467e2dc3d1fb16fbe759a1707f3edd82",
      x"861e1a822595a97202f71366a72a3886",
      x"d0de5959e75d5aa4dde824505d44212d",
      x"43586489eefe424d0ce0e918236398fc",
      x"3f58c1422eb8ad94bbfbdbc5ff7021dd",
      x"0984133c1a20a9dc777bdac6e00c9feb",
      x"3793bb6bc2e702c56f60dc66f12696cf",
      x"00cf2004bf6311e08e2314023cf6ce98",
      x"dcc3bd0d3d3bdd7c9eec9fa3795ec103",
      x"72f4a4c35c69ba460909beaa03954611",
      x"d745c917ec2647f3da7cc0a2cb803646",
      x"956998d801791174734638fff462d53b",
      x"dd6439566564747194c50ec718eb7bbb",
      x"6e2d5f55db4a381e84e66e638ea6af81",
      x"9c1dafed697cb93c20a89b11d1b345d2",
      x"a4ccf9a03b6215a421a2e06103c63ea9",
      x"cdf7162342df7e1b039fa36da5b20e8f",
      x"4275df2f25efab0b89321c9c78112e48",
      x"303adeeff1ca675735722fb6d859e047",
      x"67a95ad47b91d83c2fa5b1551058c056",
      x"be07f4ee32d6d9c763901afea74c03fd",
      x"c9072c3f66326dce2dea9acbbf715204",
      x"00a767d2d0e0b4686fdcafcff8797e28",
      x"c33798a840eb3a18ac71492132013c81",
      x"bc35c4b92c019d00109a78a3da991a4e",
      x"17e58ad81c7a0548c18951081871b2af",
      x"a1465703fda67a2e91c36445ac7dcd9c",
      x"d5f281a354d87db1cc2b7eb3c3a1f1c5",
      x"444453cbb66b6f050341e85efc4fce7f",
      x"13e60d2c839261219cea26ac23699064",
      x"0d1a6e148bac1357f07c903c5e64f4e7",
      x"02422f278683ca0c9cc7ec7732f48f46",
      x"9b16bb3faaf5aa05a9418b8b72dcc2ba",
      x"343305b12579f6ea08eea4d844025cb3",
      x"36a845cb0fe66b4ee059522862bdd12b",
      x"99364efa5f7b4022bdd930a01fbf4b04",
      x"ea08704f4051dec7475b74a475434960",
      x"472447218ffeb0622aa96cedf876eefa",
      x"a82ba271884dd96527bfedbbbc4e3cea",
      x"c9fbe12ef2e7ef724386aba4843c8cb0",
      x"bf96a0115283b432bc2b13cde9bfd0ba",
      x"05478a3cdf2fb68df93538093b955239",
      x"80ff49652f5e92f6752ba7fdcc2cfda1"
    ),
    (
      x"4e0e36136cc3c09f5843fba21efb56b7",
      x"4af7bee62cce77803255581cb15f8a2b",
      x"2c048ef5314daa5c48bd63cb239778ed",
      x"412a155637980daf24ee4ddbed0b67dd",
      x"e91c40f8d5768a5eca8e4b9625b352b4",
      x"a4e69a1502142f980617cf2af8d37e66",
      x"0e08589d1dcffcff54012b779fef9e99",
      x"7d33040f4f7e48188bb99437e436b844",
      x"7e49e66adbe92903f15a50e48d0db3a8",
      x"6a5193c4a6346771a996ba19e352ab82",
      x"7c3107c3fd982bfa43f7f2ece663d449",
      x"9eedc7015c8d7467b56d39c50150eb74",
      x"a4f7150f1c49c5ff7bdfefbabc67de7a",
      x"4b94984385a0e30c6b1d8b98fd0bd14d",
      x"c41b626577e28c3f5f61e5833687cc95",
      x"bbf6918fb0c355bb07210c2525b31f34",
      x"ed89c975bd980624ab7eb4d5c0c5098e",
      x"cc714a86637f5f39e9659a02b2ab8a1d",
      x"c3ddf372ddffd9be9b3c91fdd0afd412",
      x"789cdf69c2ca1caabbcae6d0eb4a68d0",
      x"19e335fc3aa5cbb31424db6cc8419fd4",
      x"0b438ed3ee5d0fdf7f1c39f714cf712a",
      x"a74d1f3adbf18084140aec5fd39edf84",
      x"69ff2fa71ac95f351eed3ad0275573b4",
      x"209625be6424dc61e6f60f808301ae7d",
      x"5ed20134585e2ccbd1b15f6ee57f751a",
      x"f16554e7a813d77e20d67efd86643675",
      x"d28dec643645a4c9ee1e42df44063a7a",
      x"3409e64240b1839256630666cd39ec3b",
      x"c65cb6f998ee64055e655890e310816f",
      x"152e641e14d3eee5f85d12f3173dd6ea",
      x"03b47d2c82a94d40ae3b2bd35334e875",
      x"813278f43f3f3cb2dc599966e6b6c968",
      x"5c65cd15dfd85f48b8bb39729d271294",
      x"e84215be2377fc40c0f2e19c91dea4b5",
      x"5a5cb422a35834e5353f8bfe67f8d87e",
      x"5495923cfaaa45ce56bf8c08ae7975ea",
      x"7532daa105a403abfdb67ff3db240dfe",
      x"cdd9e549245d325ee5c59584c414337f",
      x"500cc072cd6f3c0c4b0566b18bf0a5ba",
      x"1a7e5724bf835b89f0e7ff38f09cd733",
      x"923575ac39502212a88c77b2414201a0",
      x"f201b6e72d1e1a535e3ae5ce1c4f94e3",
      x"9fef4b9acaee2383b1df579e9ed86036",
      x"2e884a6b4edab626eda4654ee167fc0b",
      x"36ed89e8143fb3b13f3d90887fcb596e",
      x"72d8f0ba20027c2d3485ad77886addb9",
      x"f8fb2929008189b07e4d2344322d55a9",
      x"e03f6034e9a91715e5eadf0aa481f756",
      x"c981c0a65812903f88865514691215a4",
      x"6c27507ccc64b6cc807e44228d6face9",
      x"c6fef760eff7faa5838840deb84281e6",
      x"42b4831dccf302fb3bffc950c3da4009",
      x"c84526c7447fc2a856d96b09426fba6b",
      x"4444614788affc9c63a6fb0e00646ea1",
      x"75466f193a802d06a3609108d8e60fbe",
      x"e82de151f8b5b0cf3a0f2a5d8ac6f3ea",
      x"6da15a1beea6eb03a214b4c89b4ab910",
      x"b63df0e63aeb474a36fd39d20aa5ea11",
      x"bc5fe1f5df5d3aff594de3d46e6a09c1",
      x"54e20f3c2ed69aa42057b8730421a7d4",
      x"ffd52535956fac951f0f0cf29e5eb724",
      x"380b48602cd84d7617f396c20b02d858",
      x"cba7c6ad65cfc7e868ad4f3859b30c76",
      x"fdb3aec331db93fbc7f60d79fe13a421",
      x"521d87595207214be7cdfcf0806e0501",
      x"2dead0a84ce1ae04b36f6fa49d6bd680",
      x"cf7f1d675cc2d9215fcb169bf382d9e6",
      x"b9575151be43efef5a5494e73811ae3c",
      x"c123e038a94515769e282662301631d5",
      x"edf132121f2baea846bc5f85ba6d7dfe",
      x"786c07f8bf7938ece8d2fcf1ff3338e0",
      x"3e6cbd59759d445b4ca84f8edb72fc55",
      x"2debff18e351e030ab7e0384b3733229",
      x"4a45686e57f5b5df62668a0e84c59334"
    ),
    (
      x"56b337951e2e829cf89c0aa005fdfb84",
      x"9d70a5442be742f62805df556e36696c",
      x"e431fac2439bfada3d8dbed199b6b4ff",
      x"e389368506aa7670111dfd285afe4a5c",
      x"f0ba23b7c6c1a14b0dcc60822cf0cb87",
      x"9baa709c2328539ba6a4916fb4e0c91f",
      x"9ee60f0efa4435f8b2b68f6ddaf92799",
      x"a972a9ddb80f249690da27d6343f6491",
      x"a3f17146a78634ef18e98d1408ba2000",
      x"3ee5068eee0081856178968d160bb7df",
      x"48aa83b949aedcd68847909f4d9cd992",
      x"a9557e674709d624de84274b548d44d0",
      x"39d15aadc03bae0fcad74a43d02de246",
      x"af4c2ffd5c49ffe8c0f48ace1fcd5b85",
      x"f1592605052d3c1fc35ec34456391939",
      x"03b23a34144d2e18208adffe9fe08a04",
      x"b823942a55971c9b2fcd1eeb4ae26d3f",
      x"8b42699dc5f490196394c00d434e124e",
      x"409035d4aee93b38c4f6f13169e9b380",
      x"6147203076793fba118c456e91b3d598",
      x"33a77157a71b9f42ce79bb6fac6f5454",
      x"442d9cbe9d45647bf6baa46a58451f83",
      x"72b56dac7afe0eb623d7ca4543da8ed4",
      x"83d322ea6befc08d0512433734cb93fc",
      x"93c5cfd36fe98b115e5b28250d051873",
      x"33e914a57e5fd594ea6bad1640f6aa77",
      x"fb9213d8e1bcfe356ee3f789e3ff286c",
      x"ed9339e87c0028d7b8eeaba77ab9d811",
      x"0451362f95bb716cfae09d3d4b67b939",
      x"2400f3eb2b776e5d73634029cc738d4d",
      x"c83928e4808a43821604e53acd11bf3f",
      x"8690ea6d3d15eae85c0778f7a2200178",
      x"cd91b502fa6296abf2e5e5e9493dc4d8",
      x"739b04f0d1c32224cab4f3f06587409a",
      x"4410bb791fc422dbab253431118aabaa",
      x"177eaff71417d9c5dd983b66d3d8a64c",
      x"4e461f9173ee65a78a238b5d0dd946b3",
      x"8a7a4b05dbc010907ac8c1bc684cfb8a",
      x"df78dfab42d21dc9036c10019402c5e5",
      x"c60efaa63478c24ad660419cd5cda1e2",
      x"d378086123945a15585bdb7cd0d6019c",
      x"e43402d07fa24e54c05d08c44bf9a8e8",
      x"176342fae39c83f9525beb176b488d60",
      x"9fb058fd1a50096f808a1632f7f842a7",
      x"df543573adef123f220850b306b0f6cb",
      x"c94f3084d0487e1655cfd0b63a15cbb1",
      x"53f5639896f5eb9acd7f10d8f6bcb362",
      x"bebd7d883ff95528fac715b0578d9d45",
      x"2a77f382811909b013b2837ff27ddf19",
      x"643415536356d0d24b714d1bb92a8a3a",
      x"a2e248719ea5369c5707a004dba26792",
      x"bd7bb09c410a0f63771b2296cb5984b7",
      x"13debcfd231415f1048adf42ce5eb982",
      x"1473ce3c981e3a0fe7a28c6379f118b5",
      x"d965d9fd0242da022952044ebb38b83e",
      x"47ec9db39561e1cd5a5f66ee772d6faf",
      x"169d645e74c299093c2361795a0230ab",
      x"2155007e6b6705fbaac43c8f7e032f11",
      x"8feb9d27f2228f0b8fa191ad3a6a029b",
      x"cc8826a991db48db0542033508fbe3b0",
      x"b3caedc5268b46fdba8690005a5cd678",
      x"35e54138228f80b6d40b2185cd446f7b",
      x"5137fba76b88ab7961116387f31e5a3d",
      x"8cc586fbbd676baeb4fe3d245e826fab",
      x"03cb1dc1be4fa5ced995e85f54b62d3b",
      x"55b2373ed44d06051f85d423b5a5ef20",
      x"65767583c8c886a73fe487ae02feacf0",
      x"77e50af519adc45936316725fabf864a",
      x"987872da45f0e30069aac6e4dc30f56a",
      x"b3d19aed6e6bc8110b07151011f59288",
      x"74f0c89403358893722c10b3ab6cf52a",
      x"4d54ee1a1e5e53e92d38dbeaee3fa609",
      x"e6f1b6671c9d14b463d2cbd335444ecf",
      x"5b04b1bac70332a42bbe19bebbd44ee1",
      x"d1aa5e08afee1de8f633e6733724b24f"
    ),
    (
      x"ea6bbfec354a43a6956ab3addb60c97e",
      x"a248b9913315fd1d82df7722b212b9f0",
      x"d94b177f88de4eb5bfd2742566069b92",
      x"948191ac106208cd3fbee90a307b89cf",
      x"3ab791c8d27d1bce8b9e3476cbb5bd10",
      x"1e85e28291cc594613955bb65777a33e",
      x"a36f327974deeacf03d6e13e89283c3e",
      x"73ec71d24433b91bb1ea7bd0fc1cb4d0",
      x"67765dad0c88c43616c6208d0700d963",
      x"24fc82e708460fe13861efc330f649dc",
      x"750e822b596b7e53450ecab956903bc7",
      x"926a4c6ba97bf0a7b5848b728fa7029a",
      x"98de241e85f8d4f46e0152564b74c952",
      x"d4c7aebae8abda974b288e53ee41241c",
      x"daa9b3e0ed8bbe92641946c7630d0423",
      x"d8340587ef5d12d3804e5ed47eea4d87",
      x"1e0131068a8865dbf70d2210fbf77b06",
      x"0b1f178954640f2f64d063fb28c05722",
      x"1f43e3462687ded4146065745f037ef7",
      x"ded9b7821df51fccb0a0d898b51d90a6",
      x"6d0b2adf8fe4d8266f8c5d03c484933f",
      x"836f573683e083835b664a283eb23391",
      x"dc5241d468eaea196d4127a506cd7ce8",
      x"a15fbd15cbc48cc1d2c2a8bf9a4dd585",
      x"3b87b367156d0d540b550ac873831bbb",
      x"1a5ecae7777b25245bd0959dea5458cb",
      x"eaad195d585754bf57f9c35b4a753c34",
      x"a00ffd9552878a0d1182c6864254a0ed",
      x"4a0d375a2e6290e5d51896258142023c",
      x"fce9c198e252bc6e62b9b7061b2b21ed",
      x"50513ac4a747441ffa318d440156a6cd",
      x"e952a141151c8cefd9b925b9f27a25b3",
      x"28e3eacf7c943449f5c2a65677a33135",
      x"df0ffcd7f4130050de44784aeac5e0fa",
      x"8d59f6bb336a30b5864bdb00d4f089cd",
      x"549b56ea2a8a88740a3ed0ec7110b7e7",
      x"817c753dbf0510d92307490c59b877d5",
      x"5c380e2e4d97244aefe599b2da8bcfe6",
      x"a2e7c1f6e5ee78d1390227371a7c7da7",
      x"74cedce4546d38f6868de2bf4c2fa953",
      x"9d5f4b0b14015dc7a290351044d3df24",
      x"c9de906e4376b6e985bd10317265158c",
      x"6fb39c5f130f3e9cef6d164c32a476ff",
      x"bcf7158815247577d8dc8c69c47919d3",
      x"face43eb0589f5a64a139005c3db2742",
      x"89debf6634098091d8fa0c321d6ef7a1",
      x"b34691685b7980e27cb65b7bacc68cec",
      x"22806aafe67427b03082aafea0c92906",
      x"61b341b8fc4f9a8c5d50fc84ca928867",
      x"86020a52cf2c3e4a32261346a8d3b3cc",
      x"c1343c0294434eb6897ee4cf6962db56",
      x"034c5360c607350ae9df9a4b7cf7e17e",
      x"dba2085485d8d3ae2dce3cf35a5d71ff",
      x"18f7302be4ac78276f12b77ff82df1e8",
      x"4805b1cfb88c9d21182b90c22bba2435",
      x"35992204c9b164917c28b7cee92c391e",
      x"b237f9650b91343ccb05486f53296b2e",
      x"75d0d7ad7f6dfec429bde33834eb34e0",
      x"823064bff40276a13d857cbdd1ca898a",
      x"72e91556e87bb13f39b37a07a98c0c80",
      x"4e8a29a854141669473239bd8db9bdf4",
      x"a1d8f6850c089e06edd91177b8226508",
      x"3ffe75a5b74b6e44562703361dcfb2c9",
      x"1cb95418af95ddc39609e991bd89d591",
      x"fef3bd0b0cf30095f6e36fbedf089d33",
      x"775058a45f1290d2aa8e7e50e7cabacd",
      x"e79546c27db908c7de319726650611ff",
      x"87d1af23900d379e8228415e5019b8f6",
      x"189f73c2f3a794cde8f1c3ecec68917a",
      x"06ac11e4a94de4d30fe24f5d30a8bdce",
      x"bec9f74e4870be41a628f4e53fe98803",
      x"5bb8cca4034ba27a83139712223571d5",
      x"e1519dd834b794aa58e7fc95746df655",
      x"da0e24bbb4efe6dbed6fb1ed88d0144b",
      x"c6912538306ab0077db4c6b1aa5cd183"
    ),
    (
      x"b05c7eb8e65f32cebc88ef7a27af909b",
      x"d1162719e0f8e08d46e88d5659400301",
      x"a92ac6ea4ec2ebcbf509fc72672f66e6",
      x"84733bae92aaedf699fbd43455dc1f8b",
      x"ab71b68c7e3566f43efc7090e4fb1902",
      x"385e2b7a7590c56d7b40e9fba74246a3",
      x"90e005a066317247741716ccb8f79c41",
      x"45c78bd76bc7d02ef1728dfcfc58a311",
      x"42deff4d29c097542eb86e68faa7f7b4",
      x"d38f1cc32b62674ea4171ae26ef87da0",
      x"b5b19f6d802325ee2f73b33c96e1148a",
      x"b1f1fdf200a815ab79a947e226fccc26",
      x"4844be443d66c4dc0ec45595266b7c29",
      x"6718acd993fed8b9a4b765a43e12aac0",
      x"1375a035f25fdb128cd552cdd8ce7c88",
      x"2e8c36131775733ae5ded1d519c6c667",
      x"68ebfdfaa737ed423364258eae78d847",
      x"80a1972aad8edc7897ac26590ae0861f",
      x"1e2c02073a25084bf1552c983dad4346",
      x"8032bb694425ea66c99be19d4c871d86",
      x"ccac3ddceedb3a9b6eeec3cf993ba254",
      x"900140f2151cdf1dc4f3b9839521408c",
      x"dc6236425825d4cd95b8a90851f0ec21",
      x"d2535a7c388b30cfdea732efed94a1c3",
      x"e40de4eb0d80afdd712deaea7189c301",
      x"752edc3367ed8955b24e17311164128f",
      x"58d15eb510530f42c00e380f111cd44e",
      x"7b23fa3708b8aea3eabac6e98596cb70",
      x"8f30327421a63f60c5e5c2348ff91ae4",
      x"83b0b554eb271865b8f14f3c7f11ae34",
      x"3b961929be6544c74b3cd86cdee1c76c",
      x"8dcc278419d56dad7f1d4e7c7eeeb64c",
      x"d8d56aa216a4cb00c0f2cec7765a619b",
      x"93097e34bb695b7576a5df7cc9239b69",
      x"e3b26cbf0e8ec1278879d7fc1098748a",
      x"b713bb8ef40ffbe5d9c3381f7b821888",
      x"8bbc5f9376886d8f3628b5626d1b7c27",
      x"65e672f066036f198e9c35ba551487cf",
      x"76be8aa63c89837839d825b136ee2dfc",
      x"8f381574aac19d2f5af42699ebd9df51",
      x"7e1fea5cd801f9bf8c56cde05e5bf936",
      x"44c03874e4f03f5d9a9b0280daf93256",
      x"74ade5ee16236ffe3731419c04673106",
      x"727ec184e09b569e235d40439cf05762",
      x"4514f3064878a15e326fbdc8bb24b75d",
      x"9edb3aaf3f3b683f8f765115504d8fd5",
      x"609ab5437c33d1d8442b2d58c4d0186e",
      x"eb3783a16ba87b5ac70107cb855e97fb",
      x"1a6a50d5032a6cc6803be86f79322146",
      x"307b3f7c11fb86a7e347aef82edde396",
      x"f60db56c7a54c4505b209de8bc1e479b",
      x"96a1391dee3ff72f170f950592120372",
      x"8d758519891038a9b7859e29775c39ca",
      x"c8975e65d392d969bc7eb5143e52f7d4",
      x"a5b913e35cfdbfbb74b2236a59cf5b48",
      x"e3616058c8eef7c088cde1488eff6c8f",
      x"bd35fa7f05b9dec69d5450e204a83de5",
      x"a1620c7c58d443ff0604f6bba0287f5c",
      x"d3f0c7a94c47b5578c0a95c1f5932a71",
      x"2d28e3c4f2d96c2d8bd3a521a82177f6",
      x"9c517f4484ae8f600fde5f6ad95bc482",
      x"0d3aef0edbab78d7d4ca878e6e6c47d2",
      x"50ea6aad7e8a8f020904849e502edb1c",
      x"968a55fe5b06609bcf66afc37b5f0518",
      x"b93dfcf03a7d64ff4c332a48cb7170d3",
      x"e20aa5d2dcd849186440eecb9f313b8f",
      x"5d1cba825410dbc4612ad020012a9433",
      x"1f585bd7ea545202c6e83a743fccc60e",
      x"b932f24d70fc24edd30ccd39df95690a",
      x"777601bc91247019bf3963f7b40f86b4",
      x"fa583560833e9978673bf02a36fb5e10",
      x"fb636a1f2c41e597611d127e8959027d",
      x"cb4cc9f0d2ce657a872b1f290be86d8a",
      x"77c468f46bad95331de32619eef99a19",
      x"e8e1e755756cd4aefc822df1f1f9cdba"
    ),
    (
      x"78cc6955f2c40321af26f697c5377303",
      x"ca88b26d8e376e069a9b63c55d8256a0",
      x"cde698a58e98e938a287511239f3b1ce",
      x"b54ee944e9dd3cbd9c31e215e2ecc789",
      x"e901cc57302a299fd0cbf7c3e396b471",
      x"03791a234feec89eb78af542ec3ec421",
      x"363e7c946115612282ad051069313e93",
      x"c14f1483bf18b0f41c915aa131d298e9",
      x"a966cd4376fcf141dd5d792ee93a7da2",
      x"1ad8460bef7be26099ade8b87f35b00e",
      x"858c2270b016482b3f0a0bb45021233e",
      x"d3a4956da8f5347228e7963a06182b8d",
      x"4d382fdd82ad8d5c5762771b4ce7ef7e",
      x"a6bd26fb0219a9dc8950295d73b6ebab",
      x"78d097c50c075899aa6d9ed7177c34d2",
      x"093ace20913a333268c643efd5227180",
      x"26ed3a9dbacc91d3827bcf1d34db96d4",
      x"d8d55776956870be3281cf8726c5bd3a",
      x"eccd6b8b08a01bf4859fc7bba7baa954",
      x"ba6c435939e280e9eae5782d120f2a0f",
      x"2fbb7e62a9a9cb813da6b0d56cdbcaeb",
      x"781a9d48f1d9b73af4bf5f706ae5099d",
      x"84026e80a37f9a90001da9e0f8ed8378",
      x"6eda7e1ae1e66d00627ec8567e2d3a60",
      x"e4861080975ea85fa25532b286aa6a54",
      x"dd596bbbb640492ebcad0cfd8c3e0095",
      x"5ef4a5330dfacba02d540527140c58d6",
      x"ae19aadd16665976d19d84bd47bf29d3",
      x"46254133d7ca32d2fe4e63b73919bad4",
      x"5a300fee02209e9e4e0106e12a90f5f4",
      x"3de69f7c884b3ac35332d5e4366d3839",
      x"7ef2434a257bb04fa1acc100ad476f46",
      x"1d2cf2249c01214a693dde97aeff9ff2",
      x"bbb5e335650bdeb823b1ff089f00b27b",
      x"2c0b83d4875ea402856a114f61cf1e30",
      x"6af4f3d484fd023cdfbaf85c4e1dd01b",
      x"494480bf196ab654cae5ef36104a9119",
      x"da8604270eb00ea96bf03b3a2f260363",
      x"3afd6d209b00a0853d663ff302a00331",
      x"621e008b710b04fef498dcfb20e7f629",
      x"a253b4b6002326193d63e3a60b0d3a3e",
      x"b3a6b2bbee5197b82a04be888373273a",
      x"28d50bd43432f2969cf6ec0ab76f333c",
      x"8061b4af8565359a9e553e1113b83ae2",
      x"eb32fce73df5ced29107fcafa1363918",
      x"7c3edfcfbc9eedff8487632a4b2782b6",
      x"cf0adec390684c63fbbe65895b4f4665",
      x"227a79c555b28f466364e2c48de5bdbf",
      x"5339c2dea856286d071566e72cc47110",
      x"fc84c5dbbac14586f9217caa977199de",
      x"6d9d8627378c6f03b62b8f49fa279cbd",
      x"16efd359da865b14cb31a6a3019d634b",
      x"fb1a275aa627b5945873d454790ce29f",
      x"49febf964735f1085eb3da09e6232d24",
      x"657256c6c500b346d3b932571f3e7eac",
      x"cee897d99ed5a1d744a1a55cf0f76e33",
      x"8ac3f711ff8db368ed7236712329b30b",
      x"ce48040a2b0dba3bfdd8d7bb350d185f",
      x"9dbe53adab0bd5c780fc71a680e7b808",
      x"6cc0956b2c503982da22e0f6d65b9e43",
      x"a32b78d7fc23ec555692c06985181d37",
      x"b1fd574c01a54c16dccd901bfce0b88e",
      x"e039c24929472477020de0bf1aea5e89",
      x"97c4291c3bf0897ab92394f47894a27e",
      x"b9abfae1830c380803c133ce538f5171",
      x"ec01679e66b02f39962f1e5658ac63cb",
      x"c76cbc84780cf9d7fabd498b356a8071",
      x"9b5d9c0c8fa932312df998c2649075a0",
      x"6331962eabcfd01dce07ac773b85bb62",
      x"5e79f8190f99efc76fee42e667dc281e",
      x"f76c0920dfd29a738109b83c468c2f22",
      x"4490962c56e345db94542f24aa1f3227",
      x"d6628e6552bf205bdfc4b1d1810ad116",
      x"a753218c3b1755547ccb8b6ca1928577",
      x"6270eeda2bb3a83cdf8797acf4d4331e"
    )
  );

  constant C0 : std_logic_vector(N - 1 downto 0) := (
      x"0000000000000000000d9f6a83792fa0"
  );

  constant CONSTANTS : T_RS_MATRIX := (
      "010101011000000110101001101111010110000111001100111100010110001101000011010",
      "010110000101001011100111010000101110101000110110111001110001111111011110000",
      "111011000010011010000011011110000000100011010110100001111001100111010111111",
      "000111000100110011101100010111000100010110011011010010001000110100101000100",
      "010001011100100110101110001100010110101011111000010100100111011100010100011",
      "101100111001110011101110111111111111000010000010111101100001000000111010110",
      "101100000100010001111000001110000010110011111110000001100001100110110001110",
      "100111011110001101100111111110001101001110101010100011110100010110000110011",
      "101010111100101011101101110111011101000001111011010001101001101010101110010",
      "101001010010010001010010101110101001001010101010111001101000010111010010110",
      "000101100001111000010001100000011010100001110101100100011101110100001011100"
  );

  constant ZMATRIX : T_ZMATRIX := (
    (
      x"e1a744eddff12a7ec38075223842614f",
      x"4aa032d8005d49ce98892c73d9d21b98",
      x"048f7ea6fe2a0aaef136da047154e282",
      x"316fd41310e7c7e5c09ade69d7dc2efe",
      x"4bf11f496d63a55d6b3312645476f525",
      x"ca2c51283734fdd501636c86314f108d",
      x"0a888ae95455e2aad5aab95fa2ee0dd9",
      x"e4381ca42fbd296f3a86f8e6cf76ce7d",
      x"fa357b39bbb7d4b1ed99248dbfef1a4e",
      x"e6eb95df50336d2dd7b91179e8c04495",
      x"b3a7e4dfe2239ab6926bc0b41474a45f",
      x"5f53e45d31438675eecf736affc84e49",
      x"9985ccd9af30b166fbcad48597c41932",
      x"3b5ab98696be20d509b5f7f39f37ca59",
      x"e2625964f16ecbb7d0b916b050a1d40b",
      x"ab35dcdaf2da67372442e800fb3f5eaa",
      x"053b73762eb17750fbd1453a131657c7",
      x"b193cd987a16e4385e2a965e8c4591ed",
      x"99d8b2b982fc4718db2fe5934fbc9174",
      x"744eee531a16c078db82ff6aaaea93cc",
      x"9583b4eead8d4880d884d741093a6e5a",
      x"ffc5f20a3844ff97cbfb3adb935bb494",
      x"1b63a0e23aa925c8ee28d0cede07ced1",
      x"9a49169675fbf94bbc2f69e03b781697",
      x"75714a8afe14ef166617e1dbfb2c7465",
      x"32d6cf2272a1cc53aa07b5aad4e71a63",
      x"8fe10386980551830f99994344c3f286",
      x"38de4aec2a19a50912bcb9d2a2e40fe8",
      x"efa95f2fdd5bb4fef00cbfae975900d7",
      x"50a573153ebf76ae576f15e648510efa",
      x"229e02e54f7cef8f2193ca5a6c3fdca8",
      x"3f24cc10ae5dae4545afa9a58088d8ef",
      x"e58cc92494e8d07f22c7af507b54aa6d",
      x"d7bc8879852f74502884a42994bcfea0",
      x"b39558dc8714b24ba07b796e8c85f77c",
      x"b70fd8b2ef9d279602a1d09bc2ab4a03",
      x"bab263b7b85f6dc611d2e44260bbb0d9",
      x"d7d14924c8875db54866058132594df1",
      x"722569ee81185c87baf6acd0727cabeb",
      x"474eac14c6b640ba5f0327e03b4f21e1",
      x"e89afecabbb34d4e577be32dbb10cd2c",
      x"b47c360cf78f35d4615177e075bcaed5",
      x"1bfd4d1cd148fc9c994b1514b7f94458",
      x"2e8092c4fe65b2846fb3b514c6d6628c",
      x"7724bc4ea789d7e5e5baf8872b3aa86b",
      x"1937dfa54e4c9940921f3c5421796692",
      x"34db8057ab9cf82bd4201f4d77dfc788",
      x"28ccbc181802fcd6a04bee0bf11d1092",
      x"8370019947a81d267cf8dcd8dbe40498",
      x"c55678c0770419d7085a4db47c2e8282",
      x"ef273e4ff9afccf13c5d33c7b870e7c1",
      x"e56f68f22b4b3d7755072f3c7634e841",
      x"c3d0839a423beba0c868ae2445a00064",
      x"1502ef5810a21d3f29f50cb19a871365",
      x"cbaddb72abc93466e8195df8e2be5d46",
      x"5d2929dddeeecf48e81306aadec65d52",
      x"5ca1943cd287a8174d38acfc4be8c316",
      x"847901ef1b054de6553eed6a7c794f69",
      x"842b2f82e9bffaae19a5f1fe50b04f17",
      x"5011e94850b95937adb713e74e484eb0",
      x"d43b055f152beb2280ea1bca1590268f",
      x"40060c1b4a981341d743dd1769840799",
      x"975e5a3b184ae8b6c243df5f873209c5",
      x"a007185bc452cca227dbb215f4bc22ba",
      x"125253555245044bda38336b478b2135",
      x"af02fe1bbfd65e178495aef1acdf2cab",
      x"e409e1a6f83592efe0a0e9bde7a424a4",
      x"272da408db6f954af94ade5ee41793e9",
      x"369bc331cebda5cc16a45868497de113",
      x"c3efa04cba7dd140c1e7fafbdc1e8b8e",
      x"c9e751a6ca26f3876524a0423de00fdb",
      x"d988de06b2c89315872227d87584520b",
      x"dbaa0b3e7b49c3d0c8083c23f4c3b19f",
      x"b036e34f9f1dc42e677c3e22b91d96e7",
      x"5719802cf5c3053e782ad32fdd3aef3c"
    ),
    (
      x"252e863ecdf3195d1558503e1ff87470",
      x"13f9049d21a5ee753ace4f4ab9ccff87",
      x"8a6161b75c6c32c1179513c2d542ee1b",
      x"e4e1633908747464b8b158a64783b028",
      x"6eb54cd0fe8b2e9cee9127f3092933db",
      x"887366b9abe16f9128ba289df9ef2254",
      x"df2e59af2ca9b1dab812b34f9969fab7",
      x"05cf68c6d6d251462ae0162d5c54bcc7",
      x"5b38a874a90d50e2dc12e7499404f5f6",
      x"93464e601f0a2c6c3d7b4480857c5179",
      x"636ff7f1dd4bc9c2620042399473284e",
      x"40f7069983a6453f621611db8c4ecdca",
      x"d6ef40e755f91ef207d938791fb523a3",
      x"aaf59efd51bafd29e00d4004285b7721",
      x"9af89ae1ad95af450ac90cb258490516",
      x"d6850b979b0ed4923728f661dc310afa",
      x"c7d643db04ddf1b32d7daa1367e73932",
      x"e2d7a48c5b677461159a7c0162c90332",
      x"3b99a10bd8c53ac4d229ecb4f4218a23",
      x"5869f4a847a9df80828b1176b122c399",
      x"1a8da57f27a7f5ca823d41f0be58e873",
      x"68879c36db796b85e1483b65381f6932",
      x"b5863b15acf8f9856736bfb9100c3d93",
      x"3514c11bc6bcc9e6134c2c7c19da115d",
      x"9f86c9094f0ff35a60f7006e29ba17d9",
      x"87eae5a3ba1d49326c21c91dc9013642",
      x"4c310ffde836e805b099bbd18f06dff7",
      x"b500faee7829fba147b4908716b499a7",
      x"3b6af05ce1673ca0f6df62cda2f9606d",
      x"a552d056368a1919927d6b122eeaa74c",
      x"4460f59f7cc0cb7e644a8ba3b08f3b45",
      x"031ad3ee19d4fa107b48c0e3814f54c5",
      x"1a3b5c943a2bd6595b12320f8b104fac",
      x"d68714b0b47a586361ca5f7bb59b123c",
      x"b24aa365c6c0eeb067d23ff84d10d300",
      x"e1dcf43d303e20e9734a7610a2fd2180",
      x"7a63b3a21d27a0300a40292afff79869",
      x"ae354fb21f0efb4ed6af1bc2cee21bb8",
      x"3caff05d8e9e999b5e135f0e3be4ad23",
      x"19d2e8c3a2d76d01614af69b22e88685",
      x"761b3988f70aad175d90f0d93f511ba0",
      x"136e58a74ab6dbab45cf72c6c43a48b9",
      x"47f63c2ca12cfbaac9e2e3c150e6450e",
      x"23df74260714764ac294e39201f6409b",
      x"1b90a07d68ad18354d3aa307ad5b7d08",
      x"f161866dc55223431fc59469726004c8",
      x"a63d99dedaa540aabc41172d8c6f709b",
      x"c9260cc8481964737970a401eea022fb",
      x"84500195f5b7218f4d3b33bb38fccb14",
      x"84dcb0cf982b9148812123379a412006",
      x"c89dbe75c698d2b3e8bd83ad73a39dd0",
      x"a24cad5852e5fb37ae40137a05f7233e",
      x"a21dad88aed51b44a2221f495aa54441",
      x"9312dd81cb64c850aafa975a7fd374f2",
      x"e2f874fc0b6291436e2b59e08cade87b",
      x"388d9e9a66731e24ceb7a24a5a930a26",
      x"197cb4e9e6fa2d2f47f883b3d1cb04b7",
      x"7527ff9e15ba40d1bbca43a35d955d0c",
      x"f4035d0f8f65be5ba74cd2c8a0cbf439",
      x"ace224dafe58cdb4fa15ff289a77662f",
      x"12f9b307217b42f3cbf46e1eadc08001",
      x"3b54a1fe2a0e0e691f5bfd78fca5dca2",
      x"4a09fe4afcb4a2266c18c36b93ab169a",
      x"53c29f96981dd113b1fb7af3814f72eb",
      x"2132f5025fb0c17e5fe7a108c14b5fe7",
      x"87961a1c50001fc5071c1a404d06fad5",
      x"90b348cdd194ee1308a424d2b4a57cac",
      x"ccc840fdd007d771b61eecd5817e2753",
      x"35a2996693bf5df6bbddfb495b2481e8",
      x"46c5381f445b89673cc498552199b36c",
      x"0aa108b9e981eaa3c2178c172d2c83e4",
      x"ea5f83fc2eb7d2969cc8953073e5bf3c",
      x"2d621965cdb2fb550408ba0dfa38a835",
      x"387aaf09d63ffb8b803d9af64d4e49e1",
      x"52d47a6adbcd915cb194c97f3d73664f"
    ),
    (
      x"01d0d9b3f74e89a40cfb68f75bf14d38",
      x"6af369e8d0b56df118d241327d0f1cac",
      x"c1949aa09e89870b4153709fd3d946f4",
      x"fba8bd21f9e64b15500d42fff75df794",
      x"4e2354dd73ea97b7b0f93e45bd54a59e",
      x"eeef1e7228a05a6c78e7a260347572f0",
      x"19ec7555ecdbff2ee8fa7284dbc11766",
      x"493a63b1a51989ece54699868d99caae",
      x"cb2acad84d321ba9d5d2f9c384bce0ac",
      x"2da101f3037b839893c068192462bb32",
      x"9b025f80d01584deca2fcee10662bcf3",
      x"b8522738a2633d4ac491ecafc18eacc8",
      x"c4d16214c336507811b42b0c55de5f9b",
      x"5b9a793da12e9592ebdb04b66836d46a",
      x"628a29601d28c33d319f07947c3e85a3",
      x"a5ab13f175dfbe3b82a34f6a9b213376",
      x"bfdd8411283b9d9f8dd733b7eca33fe4",
      x"945702f15a69504412d1819f7f5b258b",
      x"b6bf58f4874ee1cfaff61d3d717abeef",
      x"c17f392d0f092ebe998d237e92485131",
      x"749a87b9fccf4b80bbf7c00367d4bed7",
      x"928ef1b827740f37595202baa434807e",
      x"7f6fff9343b55e253bfa2d5449465c34",
      x"cfcda06655636c515000b95c9c31b28b",
      x"d02d5c2faa3c00a5f6ca1a912f9eab5d",
      x"3bbe9cd29ab918a873f5fd5a4db9f287",
      x"65073b6ff7872e0aeb7369c7d440c607",
      x"41217e9b2405a6dfd4be1fa5a09b38cd",
      x"eb6d8f2590e6cd739dcc7a4fc4dbefb7",
      x"dbcb8b46c9b4ac78e1c30d08c918bb29",
      x"076e796033d4a4af62341a63188e1918",
      x"760cb43a734647ee52fede13d2eca437",
      x"a1bb9fb424246e610e966db43116586e",
      x"5d513650408bb729472fb60c4ec87720",
      x"66db6f214209e55d46e27c71b417f91e",
      x"7d93c979d3217e868e7a9648b45a2bfa",
      x"591e3772c43e724e42a40afaae9293f4",
      x"04a336add1a9b98fdf29cdafac0a4b8d",
      x"dcf479d2a4f836c819e92533a2969c31",
      x"e98f8f1083b22c677143a35aeb851c7a",
      x"f3fc99b39c69302c399eaa36b62c76ba",
      x"13766a96b01fe9bf8b33225452eac7d7",
      x"0c455e3ae4449fccaf9dfd67bcbe3522",
      x"0382de6f07bfb00822fc62a19fa18a92",
      x"b5558d6510d8d89a8bb05970e4b0d758",
      x"4a13d4f530dab89a80e6189237fb7d3c",
      x"1e8d327a735554786569620a376f8112",
      x"7120a6f70de299823b062b312a5744ce",
      x"5e837e89d3e0ccd6fe47e00b3bb5d448",
      x"d9265efb410c261c5a2f42c8bcfd38eb",
      x"296b69eee876174a3e46cca78173cc45",
      x"b85ace62d0a86c6b8eae2cfe96a10fc9",
      x"dc2014352c38f6bc96f750047dbdc505",
      x"59ef42d8f978de24dc393a44465c092c",
      x"d178cc4cbe960f491ec96d275324106c",
      x"9b562d04e72c3fe32381b2fe41f58083",
      x"cc5c2d01a8ca90f699ec67705861021b",
      x"6ae16a7f511c58b6cb530ce5338b1a32",
      x"305eb0e7aa61251e63a3533d3e4e5521",
      x"b19ece20497210a666ad64088a733f52",
      x"34e0c5e076b52f6c2659aa1c01c32166",
      x"0f69ae92b89902f0def4031d3b79d667",
      x"01512df6ecd5471821a99d714dc9aef2",
      x"ee2c082dc91eb978165dc30697da924e",
      x"75641a96d0626d8fe31e79e4a5fab448",
      x"659b9055e6fb27bea401dbaaf87b443e",
      x"cd59e76648488d8975139af71691259a",
      x"11c5187bb9d2fa9b809d06aed65dfb5a",
      x"db54c702c469612ce5f09a81adf9118d",
      x"e3a69a12d3f8616d114fb1fcb83df246",
      x"0d7319867b25666af417ecf8969f73e6",
      x"b6fd486ac71a88d1da77392904e67361",
      x"e52ccad214623c6e2d7657878fae711d",
      x"1955b98785254c843558a47fb1dbc324",
      x"8f9a36517219dc9b39458fbf59e4c95b"
    ),
    (
      x"52db02df9543a5363df9bd8757c9e7aa",
      x"4a0aed9b0bb8dd5d520ca9250a860fb6",
      x"2ef4c1be9ff9571d7852f02fcf7e00e8",
      x"20a160b7656883e402b58e9917f41c10",
      x"81cd3e85d3b17dda4046bc1a334c2987",
      x"718cbc5da20af2e0c0bbd60384e66676",
      x"9e33215f545d970d5ecff78bd2ace5cc",
      x"b62914f67c45f865cae38991e377d74f",
      x"583c3fdbdeca95605fc409b094027a04",
      x"9b4bbf1557d09676a0adb1c8b01b4682",
      x"592eca5287e120f13bdac965f1160509",
      x"3d5a16af921927371450a26e3910f151",
      x"0db01480949fd450382b2d9a80f5a444",
      x"e7a1524806d09ed504a73b17f06bcfc8",
      x"2ce7af4c7640c42d8accd974534e476e",
      x"a415aec40f53b0b0a51839b00881c7d0",
      x"9db62a5dccd3b6c5c63e9ce75fde8d68",
      x"a4a5275e0cde8327322aa1a36832a41f",
      x"4601107124a74ac41912908ef347f1d8",
      x"ad7468e01e8c5e576a7aefe0b91862f2",
      x"c70e3d25e88a5dda89663b7e296af8cd",
      x"24c01f6cce2aec441a7389cae2165390",
      x"ae114bac871ace9aef9e7b661d19d019",
      x"a52a9640cccc8162383140b74c076a72",
      x"39570ee0b3780bed8aba41cddf8bb71f",
      x"e79f42469caf7a369752503bfc8b3138",
      x"c75467f40a68070cb4017d2d18507547",
      x"22e315be834ee41451377c2f16bf6455",
      x"f910da3be720afc49dd01a2250be8fff",
      x"a040b13c00e5a8e7a1052eca5e4a28e3",
      x"5fc61a8fc844898ead5fc96690122d96",
      x"870c79710cc535cf0ff015ee1fab27a1",
      x"7755c75eb3f8fd3bc47bc2b51fe0dffd",
      x"a15dd8bd08ba2e1e063e192bd65134a5",
      x"961b311b968c1adca37486b67175a1cb",
      x"dd4027b9fb486f39d4d96f26e83dbcfb",
      x"3c28104185d43e8746ac1c4b8eba2dff",
      x"4c6ccbce4d15864e03012d85d31b9e6a",
      x"3f859720418bbf0a30627e3d78ffa584",
      x"4fb647611ca7d904319bf4a10d794d66",
      x"49c91a1ca58fdde296c3d2a3b7bf7082",
      x"4ad6bd146b43bec3a960cbf40673cd4e",
      x"8fe8364800e9efc5d8ba6eebd09af95a",
      x"4726dafa7e6b5434a948ebdbc49d4c27",
      x"f2933a4f85601a86e0c4bdcc050262a0",
      x"3d9757cb9d3d02398f62a5c6c39fe065",
      x"9e42c2568f5791175da90a1a702c8e20",
      x"7e4c5b40a60c6127ee650d78e755c7a0",
      x"c4e4fcf4391e4ee4e0306b722018a43c",
      x"ba93f90f62e3f428ffe0ab38d7307273",
      x"bd58f3ef11c468b6a768057e657b2827",
      x"3cc9841bd0bd5299b9b77b953739d1b3",
      x"712bd13117d36b6a0e6687dd99faafab",
      x"f37bc4a1fce1539d18dc2a26644fc785",
      x"e339919edf6b40c177f41f083fcf87a9",
      x"032c19186b16c4b8403879f9d5e57dda",
      x"3fa740cf6fc912312885aa7a01282921",
      x"9c7d4891b36275a86cf60cb57757eae4",
      x"20c680d8bac06ed26a0cbc32758dc82c",
      x"489dcb8f7e7221045b86219ff1170279",
      x"b8e8219e870e35fa13c93ade2740faca",
      x"da178bbdb9684e5ca83c4dfc3b4371d4",
      x"ebbdc5794da5eb5d3b4a6f696bbe1efd",
      x"5da20f9bf92eb6694a94177b458710b0",
      x"99df2e44411ccc1f577583622609881f",
      x"851bc4b62d6640fb144d079ececefe67",
      x"4127d64130133454f1ddc5e470ab9cbb",
      x"0a1380f3e1bda9b3878b2433a3412f45",
      x"9b09dd1af9d2bf0c7ad714858d0b4312",
      x"3fd1599af63e5a7bb1f4106261b53658",
      x"459fff15be041f3a93ce5e8b502b8096",
      x"5c833de847ed181d66e17be876af5697",
      x"b86bccd46e6749c7c04061d255520ca4",
      x"f72395b51ec7490308f269024e771139",
      x"2f251c9563e584f3b061bad5cbd7c605"
    ),
    (
      x"b4f8fbee3ae2b69c3bf7f7856921b8ca",
      x"f2cede24fcbf6044a7d83598208f843e",
      x"303b3de55c9cfe2391b0d9c64eab9774",
      x"4a6262b69e1c2e6f191bb397200bbf40",
      x"bf0904ce081e2af4448b7d588d7960c3",
      x"b134493a8f3ab69dccedd60a91067d31",
      x"26c22504d4ed020c07e2f644562b0469",
      x"e8d643e4803902e43116e5dbb8354ef8",
      x"b2e84e0729883a02079cd81f8755379e",
      x"64aa30209caee8ee6437ec9d5e0e3c1c",
      x"4ce13f73c603b1d94b8c5e91ab489d06",
      x"dc216ed15fc2e07c1b36cc3ae0d61f04",
      x"68c3dc570e655fdf1aa47c4d8fd325f1",
      x"c1ecc041604bfcc2044767f236b129d4",
      x"403d7a3b274704006ed1235b22eeb1c6",
      x"b25d9c82177acb54ba71e0486a7cf5f8",
      x"fd4122806c59897ef4e651c8abb34d28",
      x"bc533977a44f38fdcb2dd48f6d306732",
      x"0369f0719d69c577b12b433de9029d99",
      x"7ebb9dbca8d2b079c78d50b80515fdb2",
      x"94b1c9038be88784e60e541474190683",
      x"a3983dde7e091527f270dfe17d6e52be",
      x"a9d59855342e17e780735734aa4f8542",
      x"45fdcc7e883ceacf698c23dd4a27407f",
      x"c8c33a34d12f752498ecd9b4e40184d3",
      x"9cc0678ba1fad157d8fd33614a20fa93",
      x"9477802562a0b22a309f8a2314108955",
      x"aa6ad1fa54c315dbf5b5ea309d9f363f",
      x"d01abbc605a16316d9cc014c78eeb2c7",
      x"fe8b7aa0d6fcde9b94e23702bc9edb33",
      x"5d1b532017bf13f2e0a78bbaf6ad453a",
      x"2744ba4836f2007db716d1257a45258a",
      x"feea5a7dcafe09b473927d2761b54aba",
      x"56c231a6d4f26c391812ef78d746103b",
      x"0a0b5e8cce29eaa0b6a476e1f9b97067",
      x"6a672e4f24640b5a8ff97ab85aa66d3f",
      x"1e21fc93ce46a9f1b9a7003b2d7c8872",
      x"0f727b461f5228b20f57362958fd86ac",
      x"51a6210996c9db881f8d8f261eaf6b04",
      x"2aec1df8fa166e33d65a5ce1a9e6c31c",
      x"ea3cd5b214b7dc18463ed10e358bcf56",
      x"7d714b503d408bef3f8e78d9d3c15c44",
      x"b241307e7eceda998a2726a6a66723dd",
      x"d8cc0fc00275119eb029410545f18a65",
      x"e0a42dc5f86acca78d4862c119c258c9",
      x"b5117632d30391acec0688ddf3a8cb1b",
      x"9963fdbb89e7eda1e97ec826bc002f05",
      x"c9d1f3dbd6d1d3decba715af05cef788",
      x"8950f37855b8f8c61817fd4cf279cd40",
      x"bd489105e6521b18dac586146c5a572f",
      x"d46ecdd41e40caa8f442e6363cd63d68",
      x"3d2e14e4f231028f467775e342604193",
      x"b8eed0fa6aae0fadab72e79803bc99d3",
      x"35365fbd930c9acdb4f9a7c64da1177a",
      x"3dc48d8a46524731d8e2ace4fb470fff",
      x"f2e5144b8bf04f171e8eac53fa088027",
      x"724d53aec930c0aa2392c100a30faff8",
      x"40b80d5ab21103f096cff5bb4fa7db90",
      x"12f9fac995f2b8b81128f82bc2fc4181",
      x"5cb892330c359a96c5143c16e366ce78",
      x"ca0fd233134fb01d7f615c166560d5d9",
      x"a095cc907e7de30f035a5627fdbe6745",
      x"63b37a069a8641e1eef53d9d94b6e51e",
      x"4695b3c80f8870db8850c1d6e8c97c5d",
      x"32fdac4b2ddbf3888e86ef14f0b67259",
      x"d1fd84208442ef057c9b5b6c91b5bd24",
      x"1d76b2678284aef83a7bedeaa28df4dd",
      x"6795aa2dfcfb4d899f3cf29fc0e5d47a",
      x"e2eef6e2e7f6b30830564ae4f2a78026",
      x"97a8cf137a4ff64d2597c93735621003",
      x"f999d61ec2402a7bebea94a2e0c3a968",
      x"0328106f22ebb372f882903f561c9408",
      x"6f7a49a82b087787263936de57871ae4",
      x"fbc096dd54cd82f310d571d143cb68c6",
      x"c56d52793958fcfbe24e37197c5ba5d4"
    ),
    (
      x"6fb0f2b7c04076a3018543034e0a14aa",
      x"0c56aa21f49bd668a86500e97f6621f4",
      x"b86ef7acbf1e6a2ec7758ecfc52add0f",
      x"d4020986397f2d95e178b3fc5601c4f7",
      x"a40df98465e966d5257732cbac195d10",
      x"02dbd63306ea633a742d4d76cc6f6873",
      x"1f1847ddc0eee1d0bbc5622e94378e93",
      x"3d99bece440f7e3b0645348fb2925187",
      x"c90ffba16f137c79892e85128bcd3154",
      x"ee8c0b93a982bc0e66d53a54db5224a6",
      x"9a1de538291b56bae49eb06d4c6855a9",
      x"039e07428d0550b961d152e21cda6fba",
      x"5fbb3f9bf27bfe53ffae436dd6f1f857",
      x"7d896c3067a6ed4e53878fff4bde8f44",
      x"dfe5a2b091dd3faeb272919b5994bd95",
      x"081de2f26bdbfe029b4a58c9e8fb124e",
      x"cf32776fce4be3c0f7554fba424beef4",
      x"5aa1d2924e4bb416992164eb9fdbfc0f",
      x"1abf6e03e299849a09db5cb86748a665",
      x"19617a67dddd279418cb48e73543a3fb",
      x"0af1ffac1fefc7f3918227c2c052fd37",
      x"8030ed44475d6a8bc7523da4e8ff8f85",
      x"98df8a76a60aa4e9c349c0df22d5a6b6",
      x"3103d9846502166be35c764716b6038f",
      x"a47c602d25879deab1cbf9348eb49b87",
      x"e9d28483b62345922de09d0cdeeed743",
      x"4e5daf680e414f975c5cb375f9a17353",
      x"ac473b35df8d55d89ede73a3859e4f9d",
      x"ed13410ab5041ce6bc75b204103bc0f3",
      x"435cf4cb99147f5523fa7edf3d628ed8",
      x"f1f4d95fc595577caa181804fe22a852",
      x"4ff4b200012bb899f64ecf3f54eb7c0a",
      x"94a399e1843784b29ee202c20cfcb5d1",
      x"11c561abc1ddb114d755ac3981252c55",
      x"f102690eb5db03b93e29fa46d3bcb2ee",
      x"a7fcc48da6484c9845d216e08914e802",
      x"80c7c23b265395550999314c84811185",
      x"dc7347319ec3f869277f33d87a078766",
      x"df709d65a43dfacf600f4b9b3fbb11c7",
      x"d5a913087312f9a2fe40ac0c7246cb04",
      x"f632de62c5fd1e42ad639bb031555a4e",
      x"7db7d92a9a01b8e453719b69b24794de",
      x"430e12ae83d64a73cc76803b91aaa302",
      x"e60a5b1c9081e753322b83aac39c1125",
      x"9ab45ef7d9bf355666b01de0fdcc9b0c",
      x"12b082154ffbdcf7ead664becfce1a30",
      x"d59be01c441c90b208166be33d05e151",
      x"a785fb8a67443ff55e048a047557c2b3",
      x"c54e719318465f3a4b4fd76a6a22ee52",
      x"4d99a8e2dec319293e7fde09504334a3",
      x"e24bc0b3743907115b686eb9e06bfbd6",
      x"458194f4be4f33f92c7e1cc9c27f6f65",
      x"c9c78ad718b831dc80b62ea44ae6de88",
      x"5e77a58b0417d4ee99541ed52ac32faf",
      x"4b8842dded309b6610c3ca23ef55c931",
      x"0400fc74e326a5e97026cad8f0e55d22",
      x"d63b7e835db27cb4f1dd7ad437b80dac",
      x"74d6d4127c7d7b7a94820e7cfb2fb021",
      x"6ea27f1ba30aebec07b334ad123d0cb6",
      x"9c3f4ff559c7ada0427a2f98ae2e3a96",
      x"d37b2bdb605c8c01869ec66145fed7e5",
      x"acf89f0d01a0e393d2409a36847310ae",
      x"2a7bd68f362ea55136b4d501ced2d4ea",
      x"0931894bd379264b2d8b4028b362c527",
      x"a5319fdae60d44a0872e302960e46249",
      x"954f7174ee9c1fca4e74c1dbb823dd42",
      x"07ca3019a84614a45534c0863666cdb7",
      x"ceb2a00fe3538b4af4d7ad1fd7e9c8f4",
      x"f83abbad6ac074e0f86d215b0b338e2a",
      x"e6f1f1fd7b6b36af0105987bafc9df44",
      x"500f9de49053446d388a0d1335f3c10d",
      x"7ab041bcbc6a8a11a5e637fd208045c2",
      x"991d18abf58977b133de1f33aa430fc7",
      x"80f1d55ab4c27712e69160b7a5abd755",
      x"4eec324f5cc0464ae82d178e199b0cab"
    ),
    (
      x"3f25b36faf34a5150cce3bc70061ab81",
      x"2be6870378247a18d51c11274bdc7c8f",
      x"9f1c7cfb13e0639667e0184be721d24e",
      x"03b3b320b9a3c41ea4dcee5433e78c2a",
      x"32cf3bd291d3f46346b075806bc11749",
      x"7dc4fd85bf787631b5ec61ea9c9ea0c6",
      x"8537d22f9b9df25c913384d542ba2fca",
      x"c9f826f11d108efb7cbc5df61337a452",
      x"482f4e1071f1098694a653edf5baa7a3",
      x"c471ba47889f57f483c440bbe49e5e98",
      x"04988a676191943f4f3eba5fa07765c0",
      x"17db8412b2b0a9027fdab8457302dc5e",
      x"0b2a14bec01bf852cbf499254f00208a",
      x"39da5f8b524f546995bbb2068af0e5a8",
      x"e8e54fe7075a8d423b032979d387549a",
      x"867338b4461925791a81f7e431e9c7c0",
      x"d8e6cec6954f1d910c95f713c42b7041",
      x"ff3fbc943f6e90c205a1f52fec6b3a45",
      x"583cdda06721379f5520e887b4432280",
      x"977246b816c2e75bdc3173baa2c8f1f8",
      x"9995838a0571f5af162143ceb8da4b3d",
      x"190a45849c9a8c9f447bc786d3fd1a4c",
      x"23206d8b97fad2f482a7cc9799c3924d",
      x"dd1e747475feb8aa34263f0f4f7fb41c",
      x"4b704e726368fa523ffe2ff77c36db66",
      x"5c041e3593034c79534d72e7ff83f491",
      x"bc6adceba4cde7c30ba4854195869cc1",
      x"f7f0e668430ff90fd98d979d4d0f1fa9",
      x"c9e99c5ff2b221844cc0379a00e94e73",
      x"83aca340a0b08febfee6349d57e72635",
      x"45c55f33a604b48f3fd9d477915e2abb",
      x"ee9f36873b2e4ca548154e357373ea15",
      x"27bf0a6904816de27b81484150d32176",
      x"0fe02e57b72072452b4a2e38f5f9afb8",
      x"b75463d1addfe3d6aad2db897e3d469e",
      x"ca140533e88808b70b9650e497b81abd",
      x"e1c0bf6ee6ac3a68ca034d48e3c96449",
      x"e509b0b5f57bbf59dd92bdf0432c35f3",
      x"5268866596d6ec20bc499e3215722891",
      x"4a2d8db2a0c673764370e792a074f9e3",
      x"00dbffb3b4023ca05f9568f8b6cdb09e",
      x"e481fcc9cacb546ec875352e71ae0dfa",
      x"7d6289cdf768f49f6bab4514e333e645",
      x"f9ea665dac6b516667ba68c231eba6ea",
      x"5f795ffff2c4e768afbec05c5560d07e",
      x"1b47cbfaedd9f8a2270da5d2633e4ae8",
      x"4e94d35c4596f9689912282840551b34",
      x"118853498acec6296274c70c8dea6e1e",
      x"85ec5a82d363d0c94777b5ad34eb1bfd",
      x"5de53051a917c7b9ae45ef66609889ec",
      x"c7f56947fe68f23db4da8aa4e29d175e",
      x"8c6a2f93a9844c70fe359b0ce0bf7ccd",
      x"7e5960602e07f30c3b814ea44bf8961c",
      x"4c101541ccc8e4f307d3eb0b156c527c",
      x"e2da04bc3995a8a50aaad0c5d43d7f72",
      x"69e6db4491bb02538a0020ccf7f22f9a",
      x"77c0f082585f5c5ac3597543891ddf3b",
      x"280e2ce73e162cbd52f17dcb88aa9ff0",
      x"09ed5e7cf21362f3b3b0d5429202d002",
      x"25957e96d117982e266abd5c3b8e0cf2",
      x"8bf4680f6e5782ed11f74afb18631c16",
      x"c6bfb5a9072e6799ad73c94370a1249d",
      x"5dc2c242f41bbcf067878ae43c0e874a",
      x"9957ab77387c13d1cbf8b2c2752b0ca5",
      x"2e39b6e40ff91cae2bd8199bc56b8429",
      x"01f87fe8ae69f3194d33cd16f0f41bf0",
      x"5c2bbfc7fd11a5c1aff2b9f05f3e6aa3",
      x"a3e8cb3114d6fd650297a2eb8fd7a309",
      x"5f2e6eef3ee9a6e9c09cdf7cf5a6d378",
      x"25062e2635263d56757d5e948bfcc0aa",
      x"66fa01feb7b7303df63ce596a52d7c82",
      x"e238f9d45ae458a5a4f32c83716b0c88",
      x"0d9eef26bc9a04d897b9e932fd26954b",
      x"d84434b3538eb32cd26e509983bc09d8",
      x"a8b4970bfdea73b241d744efa93ff503"
    ),
    (
      x"bd5cf9deeb7af32408183ae57d951292",
      x"22505e1587ed252fe87a89cf11bd1c11",
      x"f30a835f58013666232a9e0a2c24de87",
      x"8b93f1d525b4f99bdce6c8e63e979e61",
      x"0e2beada4323e81cbfdc11248359f9e5",
      x"168493937df684fbb8a93d93aeb14d4c",
      x"5607c080a4612bc589e1728c17e79a4a",
      x"094c1b99e0d1510b3be4e88db41a6e67",
      x"cfc04bb398ff17d34b7b864aa526a84d",
      x"96a02b597e73f54c84701550866ef762",
      x"adb039c4cf52c68b3d16f17440f80e1d",
      x"ad736ca786f0be13425faa1ef3af9a01",
      x"a6443b5c06f1b4452f18836bd52bf0a6",
      x"8065dda628c852b8ad9e2b779e84e60d",
      x"21005db7654f5b136ba73dc3b013bb02",
      x"b7d8e3b555d144ca5b8dda059fc4c19f",
      x"b43f678ad6ccb3f694ded398a531d8b2",
      x"7f32795cbcf82389a13a701f3b99a438",
      x"8d96ec689ba1c43aaa5a0b6b9b551754",
      x"ebef129fc3139510bd291e28c8304136",
      x"c29cd47120c44d075fa5d91202b9bed8",
      x"a343b702d63320d43d611a7c84e11512",
      x"fd18c0541e6465634a8804db184ee9ec",
      x"3308054326be3baa3b8f2c4fcf38dd41",
      x"6ee548691776bbc114fa52243d4830ef",
      x"41603a2fb16b0eb61c295be3c0abb378",
      x"3135436456769098444fab9ca27bfeb2",
      x"79d16188e7c96fd72d169d4d300f4c79",
      x"0c6b6e7be5ccf318c020680c3eafbe23",
      x"f5251dcd6262c640125d4e9ab21af3ff",
      x"a0ab32b0d28adb9b38a5590249bd7fbe",
      x"58b09dfd44728f4e24d97a505f133ae8",
      x"3214ca99545789f98d41e7d06514e40f",
      x"c7db663bd0af22ae639257b2209edce3",
      x"916b237d861bcc07ca71250a99c32cc4",
      x"a2093b3ffda55a82ed5a2494ddec8ee9",
      x"80e2b60d119112da5ae62b7667c68daa",
      x"742ce80cb9f1899ed476e31e073fb983",
      x"00d770c8a1744d9792c7da72b895502c",
      x"4940d7828c9a0ca35214a63d4b07371a",
      x"cbb9a0136fb87d5786f7a03ab7ba22c7",
      x"8e27fffec7a4a773d703a0b14a225c4d",
      x"d8dad665c71ac9ce652cfcb61fae18a8",
      x"c43aba31de37b8488efd24d13c732a87",
      x"ff5406829f3868364f3cad28e9cfe13e",
      x"94a41f0bcd394e3667c8a0671ca5cfff",
      x"344319d63446900eb60a8affc96cc3a5",
      x"764a3303a5e56d5b92695ae32b206622",
      x"2301aabbb454e87fb3b42bfb5378d965",
      x"c0d173663dd2311b5eec2a3e3199b3af",
      x"af7ae7f69dbcc392e300dc2736ae68d5",
      x"4aa7cc882c031ade8e88621e70d1c964",
      x"00041095f9214b6144b70932741352dc",
      x"cb24c52034cad21afd44ff56fb66a089",
      x"c2bedde5d9bf614fdbe4d191bb5f0d82",
      x"1ff378b8a263530b2331327246764e9a",
      x"365b381000ed4ef6556308a0cfb0192d",
      x"275ca24887ba7a2ac2d2f2a2a3a4e5a7",
      x"119957864149981b33152c52cd177a20",
      x"7ca97a39dc5f8eaf0c91fccf609f5e97",
      x"4f6307657ce2fe683c4be2191c6a6803",
      x"099e00c6134c61d173355be5e59b60b0",
      x"61d3a76b78b30c4c8cb953e062869d4c",
      x"13e15f39f319f4588a9f52c860f5f2b5",
      x"ac1dd4f07c90ec70eb1ff6abb792727f",
      x"62507b25b82794a026020d1b9598d3ca",
      x"861e18cb7c696fcc108a22154b4a9797",
      x"a91d3e32d0d32dac8ec1450735ba18b2",
      x"0e00d62e10ad1921d67de99d08ee968d",
      x"7d852493fc55902e2d7386682c990338",
      x"d29c8dd0090be23753c3d7d62959faaa",
      x"4eb96835426cc0a78e0576919465e94b",
      x"f01d38ce4b56c15d87decca4928247c0",
      x"849c84107baf3bd8d09503ab2b7d1cbb",
      x"7c2482d3a0c29f30d91996b16de472e7"
    ),
    (
      x"3140defa5e83e625ada95925fb29e611",
      x"1e796051bb4b0993353175f339c31882",
      x"aa0737b0886186f3aa30812b95f8f18f",
      x"5d96f567ed10e5203ac93388e2dffb6e",
      x"2c49beab35c0a211078b7369e3f1e81b",
      x"0f16e31846a5e67e3888ec884d9fa87b",
      x"d5a9a87a042bc923d46dd1343810d40a",
      x"46e621207d3965d782e731bed0cb4716",
      x"92d0469937cf74edce68756cc5a2ed94",
      x"f3dbf91d43a0886bb1cbe1ff449ec9d0",
      x"88d3f4fe7bbe8906c600d483b55645fc",
      x"1924b482cfd8b80d123c2e06ad11d19b",
      x"d85bf82e28c2635f813c578076536048",
      x"576eb471ab81f5bf462e412b85dc9e53",
      x"6b2e79cae6c410b15ad2c9f5038bb400",
      x"e36bd4df5f187ed265598ee0ac3930c6",
      x"949ac81de82390e17cc69004c52e19de",
      x"bcdddaecc38174f6f8f1b4f4b87afeb3",
      x"3c4df25d01af4577200d51e7406b5d82",
      x"7e55f6805e72c4a3e228ec6147d48ac9",
      x"669a754a8d422610a56fe1d266fa775a",
      x"edd185d07b7a8b07c2d29c51edb3d374",
      x"d078a51b9259d1467e7fb5d2e27cbdf5",
      x"94b56b2269881202811146e4b46242d2",
      x"3d95a3977b4e20ab7f8945551d8ee2b6",
      x"031fe9a4f3df764929675d56d80d8f0f",
      x"2ccff23e11731271da6f85e95ae67aa4",
      x"984f0cd121fe064a4ce7f5deafd88725",
      x"0ddd04e7584a69a29a09aa270c3935f6",
      x"ac6c1fc58e86f225af9f5570c0171cf6",
      x"83e38cc1170031ae5bd3532dbffbb11d",
      x"5a0c3b7c2ac69526af903dd0d4ab5ff1",
      x"ce60b081a79a928cef2b726826a929e6",
      x"4e5687c10b1469e1aa8ab6ef16bc7966",
      x"0750475ca81c3bfccf055f6915056b17",
      x"977f240f3733d5d7840ed1c18af94632",
      x"0fdc4ca75cc670d90613bca6a014d1a4",
      x"d96abffc65a9a92034904878d36c67c2",
      x"3bbd102a8c8173c73a761f9d0a2d2699",
      x"becde6976f62afb90e6e4c101d2104d2",
      x"c16fcc22b19c37ceea85f452e57e0230",
      x"7f148b6a911bc59eae6db83da2967c27",
      x"e6c543be04dd59935980ce4d2b94b6d1",
      x"0b86c2ca2d549f41274dbbdb9b06d722",
      x"3a4c7b816533509d33a48d21f0673626",
      x"c45fbd634034fef4392c583c08f91b5d",
      x"92e5a7dab01336eeaac7a1cfeab1e712",
      x"11930dd46527236f299a8d4ad68c22ad",
      x"9cc91433e0f45eb316e34e3c4a46e6dd",
      x"2254242cfb231b719694f2436684b57f",
      x"45cea76b0dc7f26fa60892c1e4e5b48e",
      x"6d731c9000dc702b8c08f4945ddae21e",
      x"f6ebb914f34ba50aef5d8fd04f128381",
      x"f8b296b594bd127143ed3c5ed8e0084e",
      x"3cacf11c868401924a8a6eea207c4931",
      x"d0992eef05ca6164eebd96c0fb10b6cd",
      x"32e37b004d5f1e09c3557672f7b84e01",
      x"1678081b96ce123c705971db35bcfb0b",
      x"bd0fd8a342690ee828ffde40c37437f1",
      x"3048dc9f3b17192e0275d6f1021e1c68",
      x"3f4b99cc1828aa405a52037015af66c8",
      x"d8e34ba12cfe8f4aaeb7c0c8fc253ec7",
      x"fc24013081d6289fd2da9b26fd7f633f",
      x"06d5e5969f36044ff41e142043187da4",
      x"b6a536caf243ba18360a1fa33221ac43",
      x"9bf35bc1fc32c552c2b55fc80b60e38b",
      x"b0dc980d2234ab3720227359ed8f49f7",
      x"b8a2af5d59b738aa88a1e68439fc4787",
      x"5cc35884814c12f3b2664e4676a88918",
      x"6a9ff1ba7da58ce2cbb6b663b361d484",
      x"b3dc51238369e787606d0e3a20d122e9",
      x"1c3d49ff3e0eb02ffb208ade81c19ad3",
      x"b8364a8dd868eebd34f4691b098520a9",
      x"4b59dae91a865f38809027c8d5a1c0ff",
      x"25bc7c8e195431a3475f6d483c9e4c5d"
    ),
    (
      x"a99236e51ed18c3911ed6c97f154c1eb",
      x"bb5099283156cdbc3626f9092ac02b03",
      x"7140893b0f9d5fdd3ab14ebdf2f2ab45",
      x"e6fa6eb761a83ea264d3b7ff26611f2c",
      x"7178129abc80f664346de84868d41d10",
      x"ee593cddfeda254036ffb80c20221798",
      x"cd06b59eff345d942ed4b31cbbed3452",
      x"182d18bfd818bf9056f6dc31c09256bc",
      x"f89906671dcebeaeeb7c6873d39a7711",
      x"fe4df24d84e34a7121e9603cad8ff336",
      x"55564bccd4c9c02afc78c7acbd07a854",
      x"d5008b45753f51084cdd18d557a2341f",
      x"eee97b76a9c3afa203be4ffd5ae5f68e",
      x"683fc9dbd8fb441f761ec02258701d5b",
      x"5fb92e3196e3b1617eb4b8e1d82d21f7",
      x"93ae08f434f744e234d68963b1774b4b",
      x"86d44dd03b978083ac0711d3f78be590",
      x"66170fe119e8cb8f33756376294f0980",
      x"300e6e98c72f1d9433b79c7811e34bf6",
      x"351313ad6303cae3880780017bdd5487",
      x"d1fb4ddf730e3a4f66463aa92af22429",
      x"a4c3d45897bf5d40b9f522b085755d85",
      x"23f025734aaad09068b89095eec9c87a",
      x"b891fa62f67de892eb0f56e4ab399547",
      x"555b7b3a45900b397bf2c4c3803aec67",
      x"bde8e41fda5d6148da25b7a71625bfb8",
      x"ba15be833cc4c5c62c08d568b5b2f35f",
      x"1928314a0c74e5106aea82084bb82b29",
      x"98ab0388d8187f114294701d2d211bbf",
      x"9c6fe678c981471551cea6766814ded5",
      x"9b0d8c2156857959145fa9277b49886d",
      x"833e3bfaf3d5b19ff64d0561b61af4bd",
      x"74f5d5e241ee905185c706f9476f6763",
      x"1c1073ccc78293b3cad4bf97b7e21475",
      x"9a13f534900998355b0efba3de7c3325",
      x"7605c589de3dbeb5e0a732a76c41058a",
      x"262ccb76e713bdd3d93f3f6cd8054b1f",
      x"daf05f78823127005c623f32a21a0931",
      x"19268643f3b55c93a4d14b5069d9cfb8",
      x"a50d892f1f947c3a3389e830cde55428",
      x"1551657cef51495d60503263f528c101",
      x"db5378eb26acd916c9bcfe915ff99d28",
      x"907d4b1f466ada92a89d53febb975dd8",
      x"5a29a1835e8ba0ace924308723806ac8",
      x"f485b09012646c0b3d82bfd59758a7a4",
      x"2dd10105ac62548d572b8817b5847359",
      x"d337aec0a2e178a6be68ece93823e4bb",
      x"698b24ffa44c121ee0d568d9632dcbdd",
      x"6a4a93bcf0da0d5103defe616cf0149a",
      x"0213896bcd091cbae754cec33acb1719",
      x"280a58088be8ffaff9172fd4039ca3f0",
      x"9ef214bc38560a9589e0e2ed7d506ca8",
      x"b91f4deab2acff645859851dc3707c52",
      x"a6358977fb0dcf99d8b1209813d9b047",
      x"4b587c3ef9056442eb0eb8a72eecaa3b",
      x"59cda7bebbdfa7d1bcf7b0f4ec39f349",
      x"ffc0006492242d5d29b08231c527e23e",
      x"f5f957f8ad7c09342c27db14ed80b6c0",
      x"9c01812085e252d42c605476f2c938f2",
      x"da9d867f7d19c5a84dc5f941ce0ea822",
      x"bedaf2deb846413ce3abf2b196c74e71",
      x"41b1329b79e77ff1731db603b1dd8d09",
      x"92032d2219dd962166d08810d807cc83",
      x"4fafe0dbea66337eeb2f94fa4cc05d6d",
      x"c0a7c95f9c80839e182b6adbd9434561",
      x"67ac9c88419485b578e9d1e8703506cf",
      x"ebc226df5c7d6c0f9ae8b54ac5453d72",
      x"11c82e55b3e576ff9ad0c80ec266b73f",
      x"a7e1c876bf7c3f5053ee6416035fc2df",
      x"f1e5715b649358e1d7f547c2945e4eef",
      x"f74dd818fecc638bbf3cf7a8f64978f1",
      x"a240a9189da9457ab4d89bf04a9d580b",
      x"811cfefa10cfb3dba2f11cfeba9f965f",
      x"9ff4d381a812f66f3d2a62c78094532b",
      x"76e899b32c368f11ebc4e4dddcc2fc1a"
    )
  );

  constant ZR : T_NN_MATRIX := (
      x"4d40b94d7410784fad6f9c2ad2b81b8b",
      x"6716bc1936785366dead200d044019bb",
      x"e87fe3367b71b1da0f603bb73b4866e8",
      x"0157b6d6e1e07f6f6d534d4cf9ad1bbe",
      x"553bdb732405d4b721dfc135dfbc118b",
      x"b3ce5d195b074997e55639530c5c2009",
      x"5eadd16c3f4149493a7924758924a09f",
      x"31d9c400bf6f66cd8bc320ddb90d3b23",
      x"4a41d9b27b96a848b8271dffcd878e9e",
      x"dedf2e7d7bd6c3d419286051bfda7cbb",
      x"2970121d4b9b6ac56c80de16f18f7826",
      x"c031df95234e254f3b3ce70045081113",
      x"928ffadf9dd2aafd969925ce3634c3f7",
      x"ae58590d8196792f03bf6811eb972832",
      x"61041131337e362dce30cf60c7f6f1c2",
      x"210b697723ad081bafcfa2ee3933e1d5",
      x"a9e637a808888ac899cd11e5c6ce1be3",
      x"f23ed576a3e0cf1588d8251e9ba6930a",
      x"ea79f7db9963133bdaf3d069323630cd",
      x"107868a26e9975c3fa7eb13d65c01df7",
      x"7d273bda7be25421eac5a75db6bc3e45",
      x"0d085a62e110fe117a2623bd0eac2c72",
      x"2436aa125d087e0a4d394c39a37a976a",
      x"6c8056cba4f31b6fa887effa77a937c9",
      x"f22e772414868b24beead023686d75c9",
      x"72d04d64d64dbe23ec0f82ba11c9bcbe",
      x"90b8acc2d722421f3f6057b13bcfd907",
      x"38e8b07d9444be524cee556bc1f71209",
      x"0ab20fbdb0adf3b82e257d05d9647862",
      x"eb02a6ad00044fd70267f6633056f2c3",
      x"599bfa702654110e196d7950cec8a60b",
      x"66792215518cd10fe3a60ce8a35cd9f1",
      x"6e492b371a838589b1b721a5f42d88e1",
      x"dc699bc57a0464d629876d9750062be0",
      x"2d8e7c5d6d53d6779eba7c8af642d65b",
      x"079b0741d6097ab1f31c14bde0c38c8e",
      x"b5e05ef645e5161f5aacd9bc4d97efe2",
      x"e82eef94c60c30da8d6fd787a5afa9aa",
      x"1faa9d374d610c6c3b1de7f3c5f885fa",
      x"4d660beffeaaa894f4073cdeb63c8063",
      x"069884a09e5eaed023f11b0d57414e6a",
      x"22ba56742347c0703c38b49e88ef31ab",
      x"a82f12128305496e6007894f4df03d93",
      x"6154e3834dfb40e30b5c31e5a2cb906b",
      x"abcc227f595fa7f3c306e42d186c6b12",
      x"10aa79bc817f18fde88e46ef65a5a47f",
      x"2162a356fb4a62fe1454b24c87a63511",
      x"8e81d2159086bcf4e94417633e5f3803",
      x"08a32456e8e1fd417dd989bfabb9d0c7",
      x"36417e027095d063d9ba812220ccd40b",
      x"291fb930b5c34e44abfe20f05f0d8404",
      x"9db4a837d02b06ca9fbc750f6601bd11",
      x"ca79dcddff4d7ed81649ba89955b5321",
      x"a2b6b6afa6613175985a769701c807a7",
      x"e474b10b2f91be618972888a08281c82",
      x"d66e390dee822ada0cade384f20cee9a",
      x"a17594acc92b0d094799f618427076f2",
      x"58593273e3c6ae6c823cc7c25e408d69",
      x"90d9b8b3ee63d988e178b7a33b1c6d34",
      x"2aab4abeb8af194915a5f93123b252a4",
      x"1c1db2e64072e7c5f34e902ceea0d5d8",
      x"059ba116b1f88fa54405a615b8af60ef",
      x"5e2edb079270c6aef1703b992cbed4ca",
      x"7659ba4c4d747af77b8cb48ca142c0f0",
      x"9c21a75ac3f65b9d93544bccfd1342b5",
      x"0eccca2eca42dec1cd487065b7437193",
      x"d74a64eddc3ba1d64cc72465c6169998",
      x"8f4843a1f0ff10f7d5cde22422c0486c",
      x"c26933cf9f63e5fe1b49b2d4cd1e694a",
      x"f83c49ddb593d022a1c859d7c1696891",
      x"04a5c5e7500c6811d8b4646fe661559b",
      x"f31421cc7ea7221af29f337c5a568975",
      x"5573e415560e78b4ba72f02c477e44cc",
      x"e38af697cd88d8b345491175f23f3e26",
      x"a213aa79c0b7f466e9c6f798521b90df",
      x"aab91dbbe7ff21e29f91adde4a1fa4e7",
      x"08879fd0335a72a8c8f35a97e441f196",
      x"06a5e2c9dda64da17396b3e69279232d",
      x"59600b1c5f45c0c90d6ee5ea437d00ea",
      x"a76419735a572aa0e7dfe4ffd7ea959a",
      x"65ae6061e94dbc270b587a96e27d5d12",
      x"bd75ca326c839ee2a9f4a9a55060926e",
      x"b7c5882872ab919412e711b6763a626f",
      x"a0ccad79c43c227d294a783f8a62dd84",
      x"314fceb231c8df102f21b1741f3f649a",
      x"1d54a8efda50f1ff7590e135146c20e6",
      x"105b3b8996dc33f5d303420a347b443f",
      x"c84cbcb14995f93f798fc99f25b2cee9",
      x"ef48f257a83ce252838c4d258c03f106",
      x"53100a0860f5cbc55d4721f1f1217142",
      x"e1fde5072bb0598bdc88e5c6d492ddb3",
      x"a93fafcd5c86129fd706b63e4692192e",
      x"59cb52d3824e2daf04455f95e47cafeb",
      x"04aa5ca34f94c14e94f5fe34e4c21860",
      x"1a014f9b14bc542d4c5cb8ff7475eb2a",
      x"2ef28aec23c20a4e0bf5712897fa877c",
      x"44ddc62b2f70b2f035299b2d06ce5888",
      x"0830b9bed4f802b266150a10135b4d4b",
      x"7b9994134b9e567f3e136be567285f3d",
      x"a509de8de6aa7e000d3823d249df395f",
      x"9da7a749f1339de6b32e44c9cdcf3576",
      x"0e13d0cac923b4aec921c5269249371c",
      x"b1dcef196603927fd81f91a61fbddd96",
      x"6ce582c6ea783e71c4b077a68548767a",
      x"a08ca3001d1ae222ccb327cc96a80fbc",
      x"ed5332e34b959bd1c1e2ca2f8e4f194e",
      x"0537a6d5c14c2071a4a80913634020e2",
      x"791c7d1d72e0762dc97ad1841938f98c",
      x"f79593f3efb8fbeb572ed5159142c4dc",
      x"ca8790685f115e78c1f226381d3444a4",
      x"f104814e20959b9475d39530c9a0c3d7",
      x"cc455a0bca09589be7e355577958eece",
      x"5dfac938f8bfa9d6712fde180ffec41e",
      x"3209fb071e345740c5ed03e5959fb5d6",
      x"7c04080ac95b7189eea8c191d2c92674",
      x"fb92d2adc9b11068d34f1ab2907235eb",
      x"ea86f624bee2ef2eb307db4ea2b2862b",
      x"7522b457a6bbb19fa2facf762a539ae1",
      x"477eb6e0626ba6c3ebe6bff0096d7159",
      x"a7ddd024f8fe52013f981bf983fb6429",
      x"d61b25b61ec1e6718d31b9ffa8e5d3a2",
      x"0b0e54a2e04cfd2cbea8bae6dfc18036",
      x"986ca568e664843798e812b274bea5b8",
      x"64211eaf9bf5f9c19ae5c811f19b7e9d",
      x"9534818dd795982047c08a70de7522b2",
      x"63b34eb5ad0fcf39d7498f14b3011525",
      x"ec4b357ba6107f26e23d5d3f50b28ba7",
      x"edc136ac5d91713ff39c3742ffa78e7f"
  );

  constant RMATRIX : T_RMATRIX := (
    (
      "010111010001111110110110110110000001100110111000011100110000001111111100000",
      "001111001111100111011011011100000100101101111000011001011010000110011000111",
      "000000000100010000100010111000010101101000010100010101000101010100011010111",
      "010101101100011110111000001111111001001000111000001111011111011010000110111",
      "111010111101010000101000000100001100100111101101000000011001001011100000010",
      "101000110000000101101101100001100010100011010111001010001001101101110010001",
      "110100010011001010001011111000000010000010010001010101110000001100010001011",
      "001111001011001110001110010101000000101000111000010011010110001000111111000",
      "110000001011111100001111100001100110001111010111000000000101011000000111110",
      "001100110100101011010010101010110111101101001011000001010110101000100010010",
      "011100100101001110000110000100111111010011101101001101111100000111000001101",
      "011111001101011100001010001110100101000010110001010010000000111010100111010",
      "001000011101010001010000100011001000010000101010110010110111010000001111110",
      "001010001100001100010000100000001011010110001010010100010000011010010110100",
      "011010001011010000001101110110001110111001010000101100110111111001001100100",
      "110111010100110011001100111001111001111000110001110100001100111000110010010",
      "010001000111010000000010001000010110110011100000010000001000110100111100011",
      "101101111000011001001111011010001000011111101111011100000011110100100010101",
      "000010011110000000111011111111010001001010111111001001100000101000111000101",
      "110001111110100010111001010100100110100100010101001000101111011011110111010",
      "001010010101011100111111101000001010110010000000110011010001011001111100010",
      "011011111111011000000110011100111110110100111100111100100111001011111100110",
      "010000010011000100000111110111100011000110011100011010100000000011100000110",
      "011110111010001011100000010011000010100001001100010001101111100100110111110",
      "011011101111111011110100100111010100001010100100100101111010101000100001001",
      "101010111011110000111111100000011010001011110011111101110111001111110111001",
      "000011110111111100000010100101011010010010000001111110000110001101110010100",
      "100110011100101000100110010111101101001011110011100000101100000001011000001",
      "000100101000010001100101000100101100001101110010111011101100011111001101000",
      "000101001010011011100101101100101111000111010010101110010010101101011111110",
      "000101000110010111110100101100000101001010111001100000101100010110011100110",
      "110010011011101101001101011010010101101110101000001011100111001010000110000",
      "110100011011100111100110010110001011011101000111100011001010100000100001101",
      "001101011110011110110100010011010010110011010010000000001101001011011111111",
      "111000101010011110110100101011111001001000011000001001010101110001010110001",
      "100001101010110011100111100000001110011100111100101101001001010111000001010",
      "001100011100110100000000100101101110111000111111110000000110101111011011000",
      "001010110101101010111000100110110100011100010001111111101100110001001110001",
      "111110011111101110010000000000101111001010100100110100110001111100010110110",
      "111001011000101010010100110110000101001001110000011010011111000111111110010",
      "101100001101110010010111110101000010010111101000110111111110000010010101110",
      "010101011000111011101110011010001001101000000000100110000011101110111000101",
      "001101000001010011101101001100111110110010111001111011101000111100110001000",
      "001010001111001010100001011100111100010111010101101010111101100010010100010",
      "101000111111110110100000010011110001101110001101001010100011001101101100001",
      "110010110111111111001111111100111100101000010000111010011011100101101000101",
      "010110111111011011011000100100010010011010010010111100110110011100101101111",
      "010010011010110001101110010011111111010000110111110011010101001010110110111",
      "111101000101010000011010100111011001010000000110010010110101100010101111101",
      "011010100110101000011100110100100001010000001011010111110000000001100000111",
      "110000001110001111111000000000110100100100110100011010110010000000011111101",
      "111100101010001010101011111100110100101101100101101101111110111011101011010",
      "101101100000101111001101000010011001000000001001001110101101110001111100100"
    ),
    (
      "001111110000001100100111101000111110010010011001110010110000101100011010100",
      "100010110001111001001100001011100001010101101100110100101010011010101010010",
      "101111011000100110010001000110000111111100001101001111100110010110010111111",
      "011110000101101111111101110000111001011000100101000001011101011101001011011",
      "001101110001111001000101110011000010100101110001010100000100000011001101010",
      "111001001110100111111111100100011011010100110011111001011001010000100111101",
      "001010101101001111110011000100001111000010101111110111111010010010010100110",
      "110011111111100100010111101001111010000011100000001000101100110001100011000",
      "101110111100100110101100000010000010110000110110011111110010110101010111101",
      "010000111101001101100000111001011100010011101001001011110001000101111110100",
      "100010110110110110101100100111011101000110101011010011110001100101001111101",
      "010111000011100001011001101010010000010010000111110000101010111100010011010",
      "011111000110110100001110100010100000111100011000101100011001101101110101001",
      "000001000110110101001100101001010000111100000010111010101110010000000110110",
      "001001101000001101011000110011111000011001110001101000001010101011001010111",
      "110111101101111001101010100101000010011100000010011011010101110111000111101",
      "000111100101100101111001100010101011001010001011001101000110001101010100011",
      "010001000010010111001100001010100010100011000000111111111001111001011101000",
      "100010101101000111110001100000100010110001101000101101000100111111001101111",
      "001001111101011100100001000010010000101100111111100110111110001110101100110",
      "111000111011111010110100111011111000100010010111010100110011011010110111101",
      "001110000111001101000010000100001111111010011101111100111110100111100111011",
      "111101001011010101101100000010010001001011101111111000101001000000000001110",
      "011100001011011010000011100000100010000011110000001111101100111111010111110",
      "110011010001010010000100010110101101001111010001111111110011111011101101101",
      "100000111101000100011011010010011110110100010010111111010010001110101110011",
      "001011000101110111010001110011100011001110000111101011100000101110110001000",
      "101011111101000000001100101111001110001100001100001010000100011010010101011",
      "110010000010001000110111010001110001001011001110111101011100001001010001110",
      "000001010000000000000111010111000110001000111100000100101110000101111101010",
      "101000101011111001100111110111100111000010100110011010011011100101111010111",
      "000000011000001101111011111010111100101111101101010011000001111011011001100",
      "010110000100010001110011000011101111100101100101000010111010110111100011011",
      "001111001110000001110000001001010010100100111111110110100100100101011000111",
      "001011000001010000110110010001101111110000010110110011001110111110001101010",
      "000000101011110000000101111011010111101011001110010101110001111100111000110",
      "011001110001010110101001100001100010011010001000101010110010101111110111010",
      "011000010011011011110011101100010111100001011100010010010011001010110010100",
      "010010011101101001101000010001110010001011101100100110101111010100111011111",
      "000010110101100100110100000100110100110111101001110011011000101100111010100",
      "010000001010011111101100001110010010001111010111011111010001110001000110010",
      "001100101101111111010100010110000001001100101001111001100100100100001010110",
      "010000101011000100010010100010111111111000100010100111110011110000100100010",
      "110101110110101001011000000000110111110001011101000010001000100101110010011",
      "101001111111000111101111010010000000010110101000000111001011011110111001000",
      "000101101110100100010000101100100111100101001011111111101000100110101111100",
      "101000101000111011001110011000111111010011111001010011011100110101001111011",
      "010010010101110110000111001000100101001111101010011000111110111011001011100",
      "101001100100000100100010011110001010000001011111101001110111100000100100011",
      "001001110010110010101100001100100110100010111101000100011110110111011110100",
      "011111100001101000000101011010100110110110011101001010001011111001111001101",
      "100010001001111101110100010011110000010110110000111101010100001000100011110",
      "001001010110001111111000111110011011010010000110001101001000001111010010010"
    ),
    (
      "111101110100001011100000111010110000010101010111100001110011111110100111101",
      "010100000011010011011000011110101001110111010000001101011000100011010000101",
      "110100011010001101001000111000001011011010000001111001111010100101100000001",
      "000101110011001010101101111110000010110011110010001111001110110001010000001",
      "011000101100010010010111011001110100110101001010000100010100000111101010100",
      "101111010010100110001010010111001001110111010111110011011111010010000000010",
      "010101111010110000011011100101001111100010000011110000110100111001111011011",
      "110010100011100100001001001101000101000011101011100010011100111111110011110",
      "100000110001100110010001010101000111011100111000101110110101111100010110001",
      "010100110111000100100000100101110001001110011000010000001010011100011011110",
      "110110000110100010000110100110100100010101111010100011000100001101010011101",
      "101111010100010000111000110011000010101111000011010100001100110010000110011",
      "100000010011010001110111110111001011010100110110110101101101111100001011110",
      "111010010000001101110111010000101010101011000101011111010000000100110011101",
      "110000110110100101010111101001101000000001010001101001101011111111111110011",
      "010100101010100111000101100111111000000011110110101101100000011100000101010",
      "010100000001100011000101011100100100010110110000110010001100001110011111111",
      "001110101110000100110100000000001111101100000110111011001010010000000111110",
      "111010101000011010001110010111000110110010100011100001001000111011000111101",
      "111110111001001100110110111001001001101001010101000000011110101000010101110",
      "011011001111110000110000010001111010011110001001110001001101101110000011100",
      "100100011010000001101101101111111110111101011000001100101111000111111111000",
      "101001110011001101001000010000101101000001101011100010001000101011001100010",
      "011000000010010110001111011111010100010100000010011101100111001011010000000",
      "100000111010110111011100000001100000010011110011011000000111001011001110100",
      "011110010011000010101110101000111010111101000011100111011100001110000001001",
      "110110100010111010001001001001010001001111000011001111011101100111101101001",
      "000110111011010000001101111111000001110101000001011110111010101011001010100",
      "101101000110111110000001101100001001101100101111010110110101100100000110011",
      "100011111000011001011010001010001111100110110011101011011000000100010000101",
      "101110000001110111010101110001001011011100111000100001100011110000100110110",
      "110001001001100010101111101000100111111000110011010111101010011000101100111",
      "000111000110100110011101111001000001011110000010111010001111110100101011111",
      "100111100010001000101000010011110010010111000101010110100011110101000000110",
      "000011111110100100110001011111100001011100001011110011001000010011111101101",
      "101011011010101101010101101101100110111001010001001110001101001000111111111",
      "000000110100010110001111111011101101011010100001000111001101111000111010110",
      "000111100011100100101010001101101110001000110100010011110010100011011000000",
      "001110101111011100010011001110110111011110010000111001010011001111111110001",
      "001001101110001110101100001111000001100110101101100001000000010100111111010",
      "111011110101010001111011111011000101011100001010100000000001100001010001000",
      "011000001011000011000101001111100111001011000000110110001000000011001010011",
      "100001110000100100111001011010101010101011010011001111001011110001011011111",
      "111011001011111110100101011110011001010100010110100001100100011001001000100",
      "000110011111011100111111010111010011010001001101001111101101110100011111101",
      "110111101011011101000100101101100010100001100001100011011110001100110011000",
      "001001001001011111000011001010011110010111111110011110000001000000110110101",
      "000100011001010010110001001100000101110001010001111001100111000101101000000",
      "000000000111101101001001000110011001000110010001101000110011111010101000000",
      "010011100100110011011110101000111111110110010010100101110011101001001111111",
      "101101001111011000111001110101101000001110011001110111010101011100000101010",
      "100111001101100110111011100010000101011101100100000011010001101111001011111",
      "001001010111100011000000100110100110111110001000010100100110011100111011111"
    ),
    (
      "110100111101000100110101000010100000001011100010110011001011100101101001011",
      "011110100100101100011000101110111010010001111111001011000110010111101111001",
      "010000001011110110010010111101110001100100000111111111011111010101100111110",
      "011010001000100010101001100100101111110011000110011001101001001111101010110",
      "100110001110011000000010001111000101010101000010100001010010000101101101100",
      "111111000100101100100101101001100100111011101101100010000100001011001000110",
      "011011010000101011011001001011010000100100011100000010010000001100100000011",
      "100100000111001010110111110100100001000110010011110010100100010110101111111",
      "110101001011000110010111011101101000101000010011111010001010011101000011110",
      "001000010111100101001010111001101100110100011010100111110001000110111101111",
      "111000010011111000101011111000001000110000000011011011000010001000000110100",
      "011110010110001010011011001100011111101100110111111100011001001111001101111",
      "110101111011100111100100001111101100101110001111111110111101010111110001000",
      "101101011011111100010110101101101010010100101100010011010000010000000110100",
      "000101100110101111001111000100011010010111010100011001000001011101110101011",
      "001110101010011000110010100110000101011111001111010010111100101000101000100",
      "011110001010010000100111110101111011001010011101000010001111111010111011000",
      "001001110000011000101011101110000100101111011010001011001011110001001010111",
      "000010011101000101010010011110111011010011110010011110111110110001001110110",
      "011001000010101001001010010101110000011111110010110000101111100100010011101",
      "001111101110111100011100111111000101010001011010101100011001010010111010010",
      "101101101100101101100110001101100100101100000110011001010101101110100100011",
      "100010111100011001011000000111011000010010100010101100001110001000100110010",
      "100011100001010010011110010100010011001001100101010010000000111100010000111",
      "111110010010110110110000000000000001100110101000011111011110110010100110111",
      "110110010001110010111000011111011010000110010110111111000010011101001001100",
      "111000001010000010100101101010001110000101100101011111001000011010001110101",
      "001000110100111100100110110110000100111010111011010101001101100111110001101",
      "100000001110100101010100011100000101011100111000110110101001101101000111010",
      "000011001000101001101100101011011010111100011110000000000111000011000110000",
      "101100010111111000111010100101111000000111001010110000011100111100000101110",
      "100001010000010110010111101110111100011111000111011010001011111010001001010",
      "101011101010001001010000000001001110011001101011100000100111100110101011010",
      "001101000100011111111100000001111011101001101111001011001111000101110100001",
      "000100111100101110110101111001100100110111001111111111100010111100110111101",
      "100101101011100010010011001101010010110100100000010101001101101001010111101",
      "001110111100100000110010110101100111101111011110001010011011011111101010111",
      "111001010000101010101011110000001001100111110100101000001001000011100111010",
      "101011101010010110011100001001111010110100100001101100010000111010011001100",
      "000101101011100101010010010011101010001101100110101111000010001101110001101",
      "011110110110111000101110110011000110101100110010010110000100010011101000110",
      "010010000001010010010111110111010101011110111001110011101111111001101100000",
      "011111001101101110100000010001111001010101111110001101001011111101011001001",
      "011111000001110001001100111001001100010001001010010111110010010001100000101",
      "100101001111001001111000000000011001001001100101001110100100001001001100101",
      "001010010001010110111000000011000100110011001001001011110010000111101010101",
      "101110001000010010010000001111100100000011100011010111101111100010001100100",
      "100001011100011101101110010100001011100111101110100011001000011111010010110",
      "101111100100111011010001101111101000111010011101010110110001100100100010010",
      "110101000000110010010001011101000000011101101111111011000100001010111001001",
      "001011100111011100011011000111011011100101001001010001000111111001111010010",
      "111100100000111110110101011100110001001011011000101111110001101100100110100",
      "001010010100110111010010111111101100111100001011000010000000011111110100101"
    ),
    (
      "001101010000111011101110011101010110011000001111111000100010100101111111110",
      "100101010000000000001101111010010111010000011011100001000000111001001110000",
      "100101000001111110111101100100100111100001010011011111011111011100111100000",
      "101101100001011101101101111110100100100001001010111011101011011000111001101",
      "110110110011100110001111111100011110111010010000010010010111101101111000101",
      "101010010100100100000011011001010000010110101001001100101010000001010100011",
      "010001010101110010100000100001100100000100001001100001001001010010111011001",
      "010010111011011010111001001001001100010001000101101110111110011011000011011",
      "000110011001110111110101000101111010110011100111011110000100010001010010101",
      "000110011001000101010111011100000011010110000001010110111111010010111111010",
      "011000010101011010001111001110101010110000100010101101111001110011000111100",
      "110000100010110000001011111100000100010010010101000000010001110001001111110",
      "000010010010110011110100010111001001000111000100101110010110011111010100110",
      "001001011010100000011101101100101000110111101110111011001001011101000110110",
      "100011100001100000011111001011100011111000001100111001100010000101001000100",
      "111011111010011111010110101100111100000001000110100110011100101001110001001",
      "101000010101100110100011010101111101110010001001110000111000001111001100011",
      "111001011000010101101111111010001110011010101111000010001110000101111000111",
      "111111011000001111001001011001001101011000111101101000011100011101010100000",
      "000100101101111111100101010011000111101000001011111001111000001010001000100",
      "011000011110110000000010000011100001000000010011100111110010110101011010100",
      "111010111001010001110111110011010000000000111100010110111011000110010011011",
      "101110000101100001010111001011000000011000111000101101000110101000111001001",
      "100000110011111001010001110000100001000110100011010110110010101111010111010",
      "100111111110100100000100110011000100100011011010001101110100111100111101101",
      "101010101101110100000010111110100010001010011001111100010000001111000100001",
      "010011010100000000101000110101000100011110111110100001101001110100101011010",
      "101000010010101000101100111000011111011100001111010100001110101010110011100",
      "000111011100101101100110001100010111111110101001100111100000101011011100000",
      "010110011110001010011010101100110011111000001111100111100010011100110110001",
      "110011011101011000010100100000000100111011100111010111010100001001101011110",
      "110000001010111011110101011100110111011001001110101101011001101101000011000",
      "101101100101011100101101000101101100000100000000100101101100111100001101000",
      "100110001011011000000011111100111000011010011111100010010011000100100110110",
      "110111000011111101001101011011000110101111011111110010000111101110000110010",
      "010011010100110110111001100010000011101000100100000111000010110010110010101",
      "001010110010101001000111011111110001110100010010011100011001010011101101101",
      "110110110101110010000100010010100100100000111001010101110100101001000010011",
      "101010010110101000011001100100000111001011100001100000100111101110110111001",
      "100011111110001101100111001010101011101101000110111001100010011110001111111",
      "010011101111000001110110100101111111011101010010111001010100000100100100001",
      "010111001101011101111010001010010110001100111001100000000100110000001100000",
      "011111100000011010100101010001001011011001000000101000101111001001110110111",
      "001100000010111001000001110011101101011100000101101111011100100000111001001",
      "011100001110011010110000010001011010000000100101011001110000011010111101111",
      "101010000001001101110000001010001111111000000000101000011111000000010101000",
      "011001110000000011101100100010100010001111110011111001011110101011000001110",
      "101000111111001010010101011010000010100100100010101110100110000011011010110",
      "001011100011111001110011001110110110010000010010100100100011101001100001101",
      "000101111011100001010011110001000011111101001110000010100001000010111000101",
      "000100100100100001110100001101101100100010110000001101010011000011101011000",
      "110010011100011111000110111010000100111001110011001101010000011000011101000",
      "011111011111001001110010001010110010010101101101100100000111010001001000000"
    ),
    (
      "100011010110111000100000011011101110111111011101000111111111000000111010110",
      "111000111110110110100110111000001101001001000100100101100100111010111010111",
      "010110000110100010010010000000000010010111100110000011110010001111110110001",
      "011110111011011011100001010011001101100010101100101111000010100101100111100",
      "011001110100001001001010101000111000101101000110010000011010000000100011001",
      "111000101011000100100000011100011100110111100110100111100101000000001000011",
      "011010101100101100011010011011001000111101001011010101101000001100000011101",
      "111010100110000110011000001111001101011111001101100000000000101000000111001",
      "001001010101101011000000101011101101110111100111010001111010101010111010000",
      "110000100101000011110111111111001110001001101010101000100111000100010000011",
      "001110011100000001110011111001010100111001111110001101101110111000111111010",
      "100011010110010000100111011110111010010110000001010010001011010110000100111",
      "111110111000110110000111011011100011100000100001110100010010110101101000001",
      "101100101111001001101000110011000011111100100000001010101100000010000001110",
      "010011110110100100101011111011001011101011110100011110111110010110011101000",
      "010001100000001000100111111000111100110000110100111111111110111000001100100",
      "000101001010110011110011000011011111111010001010010000010100100011000110001",
      "000000111000010010001101001111100011100110010100111111111110101110001110011",
      "000111010100001011000111000110010000100011001000110111110001111110000101011",
      "010010000001111110010011110001110110000101110110011110111110111010101010011",
      "000010010010111111100010110100110110101000101100000000111110010111011010100",
      "000111011110100101101011101100010100010000010011000101011111100011100011001",
      "000011101110000000000011010001010000010110010110110110110101001011110100010",
      "100111100110001000000111110110000000010001010100010011110100010010101110100",
      "000111110111010010010111001110001100100110000110111001011010100100100010111",
      "100111100100111010111001000000001100001011001000100101000010000101001010100",
      "001111101010111100100010001100001100010010110111111111100000110010101100000",
      "100100010001100010010011111111100010101101000010110010000001010000010010010",
      "001011110110100100110110001111001011101111101010101100100000101001011101111",
      "111110010100011100110010100110111000001111001000000010001101010110100000111",
      "100111010101001011111000100100100011001101101000100011011011101111110001010",
      "010110111110111100110000100000110111001110001110100110100001111111101111001",
      "011001011111100011101001001010011101100000101110101001111110111101110101111",
      "011000001111111101111110111000111110010011010000001000010110111000100110110",
      "011010010001011000101010110011010100101111111100100001100000101010110010111",
      "010100000110010001000000000000000100110110001111100100101010000001111000111",
      "100101001001011101111001110000100010100000110001011111010111011000000011100",
      "010010010100110110110111010011101011001001100011011010110100101011000100001",
      "110101101010011100000100111001000000010100111011100001001000101000010101001",
      "001010110011110100100001110101001011011011001001001011011101110110110111000",
      "011000100000101100111010111000011001110010010110111001101010101001111011111",
      "101110110101001111111100001111110110110111000001111000111100000000010010010",
      "010001111100011110100010011010011111010011000010110111001101111110111011010",
      "111001101010011000001000100101101101111011111000101100110111011101111010010",
      "111010100010011000000111110001111100111000111111011010100101010000011101000",
      "011100011110010100100001000100010000011001011110111101010101111111111111011",
      "100100110001001001111101000001110110110111100111010011010001000110100111001",
      "011111001000110110011100001011110101101110101111001001101011011000011101000",
      "101111110001110101101011011001000000110011110110000110110010011110000100100",
      "011100011010101001011001010000101110010100100000011100100100010010111011110",
      "011110001000011101000110000111001111010011110011101010101100011010110010110",
      "100001001101001000100001011100001011100010100011001100100000010000001100000",
      "010010111101110111100101110110110000010011100000000000110000110100101110000"
    ),
    (
      "000100111100011111000011111001001100111001111010000111100111110101010000011",
      "101011010111111000101111101010010001001111000110110011100011100111100111010",
      "000011011001100011010010011000001011110101011100100001100100010011001111001",
      "010011110010111000110100000000111101110100000110000000010010011010001001000",
      "111000101000001011001011101101111110111101001100101001100111001001100100001",
      "011100111010100110010110011000011111001001011010001110000010110100011101010",
      "011100011001000101000111101010000011010011010010001100000000101010111010001",
      "110011110001111000010011100100010100100010110110000001011001000100000001000",
      "011110001010110010000010010101110000001111011010111000101101001100101000011",
      "110101011101010001001011110100111001110010010100110011111101010011011111111",
      "001101100111011001011101111000111011110011100010110000111000111101001000001",
      "000001001100011100000110111100111011001100000011001100010010011100101111010",
      "000110010011111001101000111000001011110010010110011111000001110011101110011",
      "100001011101101100010111010110100010110000010111011110000011011100010011000",
      "110100101000011011100010000110100100000100010100111111101000101100001001110",
      "000110010010100111001000011001111000101100000101001010001010101000010110110",
      "001100010111000110111011001011000011100110000011001000011000001000011010111",
      "110011001000100111110000010010100000010100011001110001111111100110111110000",
      "101101111011100111011101010110010110101111001111011011110100000010010010010",
      "011110100100100101000001110000110101010000001000101011001111101110111000101",
      "110110001011101111110000111100110111011001010101011000010000101001011000100",
      "111001100111101010101111110011011001000100000110011101001100010000001100111",
      "100010010010001101110000101110101100010001010100111001010011101100001111101",
      "101011110101100101011100100100110111000101000110010110010011111100001111101",
      "001000010111111001010001000111010111001001001010010010101001000100000110011",
      "000110101011110110001000000101010111010011001011111110110000111010001000011",
      "111100101001111111101100100111111100100011011100010010111111110101110011010",
      "100110001100011111110000000010010100100001110100100111010010001001111111001",
      "110101101001000000010011011010110000010110110001110010110101011011110110111",
      "111110101001100101011000000010010001111001011011011101001110011010011000010",
      "000100110000011100111110001010011001100011010001110101101001010101000111010",
      "111001011000110011101110010010110010100111011100010010001010101100100011001",
      "100001000010111111111010010111010111111110111011110011010111111100011001110",
      "111001011101011010101000100010000011010011010110000101100111101111100111110",
      "001011111011011010110000010101111011110100111111010000100011001100101000111",
      "100110011011000000001110011101101100000010111101011111111101110011100000101",
      "111011101001110110010000100110101001111001000010011101001111000011101110001",
      "101100010000111001000101001001011110100111011110010111011111101100100010100",
      "100111010101010011001100000010110101110111100011111100011001101001100000010",
      "110110111110110001010000011000110101010000011111100101111001001011111000110",
      "011000110100100010011010011000110000011101100100111110101010000100110100110",
      "010000111100010000001100110110111001100101111001000110011011111111100000001",
      "000010110010000010010110111000010001101111011000111111111110110000101100111",
      "100101000000100100111000001111000111000011010010001110011000010101101100100",
      "000110111000100000111010110001101100000010000001000101101011000001011010101",
      "001101111010010100101111010011100100101011101000011101100011100101110110010",
      "111010011101000011111101100100100001101101110001100010011101100111011010010",
      "101101100110001110110000010101001100000110100110101011110001101101101100100",
      "011101111110100101110101111011011101101100011101110110010111010100100011100",
      "010001110111101111001110011110110101101111100101010011010111110111101010101",
      "110000001111101100011100110110011100110010000101010001110010111001101011001",
      "000010001100100010010111110100100000000110011101010010001100100110111100101",
      "110110010011010111111000110000011100000100100011000110100010110001010000111"
    ),
    (
      "000011010000010010010001110001100000010011110001011010010110011010101101000",
      "011110001010001110000111001101101110101101101110111001110100100000010001100",
      "001111000111001010100000000000100001000011011111101000010101010000011000000",
      "101001111101100001101100000010011011110001101000001111000101100111101100000",
      "111100101000110010110011000110010111011011100010001100110010100101100010100",
      "010100000000000000110100100011111001110100011100010100000111011110101001011",
      "101101110000010011000001110100001110001110010100100110010000001001001110010",
      "000101000101110000000100001011011010011101001011110110011101000001101111110",
      "100101000000110010000010100101111010010000111100000010111010011111111100001",
      "000100110100100111100101011000011010110011000111101001001101011100001101011",
      "001110010000010010000110001110101000011100111010000010000001100010011001011",
      "111010100101011101111100000010010100010111110111110001100010011000011111001",
      "000111001100000110110001100111100010011100101111101010001011101101001010010",
      "011000101111001010101011011000110011110001011101011010111000011101001000100",
      "000100001010000111011110001011000101100101110100010011001111000100010111110",
      "100000001001000110111100111101101110100110011001011100111111011110100000010",
      "010000111000000001101110000111001101111111100111101111110110011110100000110",
      "111111010000011001010111010000111000100010011011110011001100100000010010010",
      "010100110010011111101001000000011111111101010011100111111001010110000110011",
      "001011001100111000001101011111010110010100101011011000110110000111010011000",
      "101101001010100101111011011000111000001011011101111100001000001110001011011",
      "010010010000000100110101011011011011011100010111100001000110111101100101100",
      "101110111101100000111000110011011000011100111110000000111001010001111100111",
      "101011001111001010001100001011100100111010011011010001001100000000001101101",
      "011010011001010010000010101010111011111000010010111101111011010011000101001",
      "010101101001110100111111001000101001100101000001101010101110100011111111110",
      "011111001101011110001010011001110101101110010011010111111100100011011011001",
      "110100000101000001100101000110101100100001110000111111001100111101010101110",
      "011101100000011111110111111111111100010111001001100001001101110110000010010",
      "010000101111110000011101100111101111111101101000000100101001011100000001000",
      "001111100010000110011000101110001110010000001000110111000000001100111110010",
      "111011100101111001111111101110010100111011010000001010001011011011100000011",
      "001010110111111110010010111111000110000110001111100010100100011011011101101",
      "110100110000001100000111110010000110101111000000000000101111101101000011101",
      "100010100000000110001100001001010111010100101110110001101011011010110011110",
      "111001010000111010001110100000111111101000001111011001100001111111110000010",
      "101100001111001001011111110000101101011000010011010111000110011111001010110",
      "110011111110111000110001001001010000010000101000000010001111100110101110101",
      "010001010001110100000001000111101011010100000101010111110000100110010011001",
      "110000100010110111010110110000000010100010101101011011001001011110110111001",
      "011001001010100100010000110010100011101100111101111110111001100000110011001",
      "110110111001001000010110101100001110101001110011011011101100011111100010000",
      "010100110001110000001001010001001100100000000111110110101010100001011100010",
      "000001101110011100111110010000110010010111101000010001111011100111000101111",
      "100000011111101001100110000011010101101110011010100011110010110111101100101",
      "000111111011111001010111110111011001100010110001010010101100111111100000111",
      "100100100001000100011100100011111111101110000011101100011101010100001100000",
      "111011001100010000100000110000110010000100000100110111111110110101111101101",
      "110001100011101010000001000110000001001010000101000100010010101011110011101",
      "101011111001101110101001100111010000001110010010010011010000010001000010101",
      "010000110001011111011000101101000010000100110110100010011110110110001010101",
      "011011100001011111110100011010111000010001101100001101011010010100110011100",
      "101001110000001100111111011101000100010100000011011010100101000101001100111"
    ),
    (
      "111101011010101000100000101110111101111011100100100011110110000100010110010",
      "111001111100000100000000100100000000101111111111001010100011001101001010110",
      "110001001010000010111111000010101010110001100111100111001100100100111111100",
      "010101011011111010110001101011111101001111001011010111010001001001000011110",
      "101011011011110010101011000100010100111110111011001100001000000110110101111",
      "101011101110011100001001010000001110101101110100110011110100000100001100100",
      "010110010011010100101001101110000011110111011010001111010111001110010010110",
      "010110011110001101101101100001011001010111110001000100000100000111111000110",
      "000001010000101110110001110001010111101110001110111000111001110011100101101",
      "000001111010011100000001111101101110101001011101011101001110100000110110010",
      "100010100001011010110100001110001000101100011111001110010111010000011111001",
      "101000000010101001100001111010110101101000111101000100111000111111000000110",
      "101111101011101111000110000100111011010100001110011010000000001010010011010",
      "010001011010000101100011001001101001000011101101110100100001011100101111001",
      "001100001010110111001110010010101110100101110100111011010011110100100111101",
      "101010001011001100000111100111111101010011101011000101011111101101101110101",
      "101011100011110110100101001010101110111011001111110001110011101010000100101",
      "111011111000010011101100110010001000011110110111100000011111001010111000000",
      "100101011001100101110010101100000110001011010011100110011100100001000110100",
      "011010101011101000101101100111011101010011001011010100011110111111000111100",
      "001111000011101101110111011100110010101100010001010100001001101011000110001",
      "011101100101000100110100000111000110111110101001010110101110110010100110101",
      "101000110001001111010000111111000010001011110100001100110000000010101100010",
      "101011111111111001100011111010101011001100110101000100010101100011000111110",
      "100101001100010000100100010100011101100110110001001011110001001001111011001",
      "110110001010110111110110100001000001110000110000010000101000110110111111110",
      "100101110001110011100010010101011001111101111111000010110001100111100111010",
      "011100001110000011000111111101100010010011010010011110001000010001110011101",
      "100100001010001000100111011110010110100010010001011010011101010100110100010",
      "000110000000001110110010011001010011010101101000000110010110001000010111001",
      "100010010110101000101010000111010110010000110111111100100111111101000111111",
      "001111100111100000000110100000000100001010110110111100110001010110110101110",
      "101101011010111001110000101101101001110010000000010011000011001101001101011",
      "001101001111111110100011100100100100010110011000110110001010101000011100011",
      "001010011000001011110101000000110011010001111101110010110001000001101011001",
      "101001011100010011000001000101100100110001001010011000000010111101010100101",
      "100011010000111000100100010111110110101000101110101011010011000010111001110",
      "100001011111100000001001111100001001100111100111101001110010001001010111110",
      "011010010000000011011010001000110110001100111100100100110100101010101010011",
      "011101111001100110000011101111011111010101000100010100001011011101010001000",
      "000011100011101010001010011111111010100100110001001111011110101001010101011",
      "101001011010101111001101100110001110110101110110110011011001010011000010101",
      "011000000011110110000010001100110111001111011101110000100001100111100111110",
      "010110000100111101110001111110010111111110100000000111011101110110100101001",
      "001000111110001101110110001001010011011111011111100100000110000010001100011",
      "001000001010110001111100110000000111000100011110000010010100110001011011000",
      "111111000111010101111110011010101011000110010101110101001110010110100010110",
      "010001011111011011001101110000110111101101101110110110010100011010001111001",
      "110001100110000011100111101011111011001011001100011000110111001000101100011",
      "111110000110001100101011001001000110100011110111100101011001000011000110110",
      "001101000000000100000000110010010100001101111000010000101110011001011100000",
      "010100000110011110110000011111011101111101000110000111101101010110111000100",
      "100110010000110110000100101001000101101111000001101111001010101000111111000"
    ),
    (
      "001011010101101111001001001111011011010000010100111001011110000011011011110",
      "011110010000101010001001001000100111101001000111100101100110100000100000111",
      "111101010111101001110101010010000111000010010100111101111010011010101110000",
      "100100111010000101001110110010100000111000011010011001011110000110100001100",
      "011010100011100100000100111001111001001111100100101000010110000101010101000",
      "010100000010010011101110100001001110100100110100101011010111000101010001100",
      "101010111001000100110101101111101110100011001000110111001000111000010101001",
      "011001101011001011111010101000110001011100010000100001000000110110000110011",
      "000010001110111100100101111011011000110001101011100101000001001111111011111",
      "000001101111101001010111100011100010111111000101101011100001010000010100100",
      "010110000011110100111001010000010010011010111000100100010000111101110011110",
      "010110100100011101111000111010001011101111000001101101110000111000101010001",
      "100011100000011000101110000001110011101110110101111000001001101110111110111",
      "000001111101011001110101001001101001110101100000100011001011010111010010001",
      "101010010000001001000000010011101101101011000101001101111011110100010001101",
      "010000110101100000001001010100110010100101000001001001001001100100110110110",
      "101111000000101000010010100001110100110000101011111111011100010110100110000",
      "010011101110000111001011000011001110011000101010011111100111110000100100010",
      "110111010101000110001011011011111000010000010101110011101000110000110101010",
      "001000111101111100011100101000001111110000011100101101101011011000111001100",
      "101001101000010110100000010101000100011100100001101100101100100111111010010",
      "110100010011011111000110100010011001101100111110100101011101110110010110111",
      "110100000001001011010001111000011000111001101101000000011010110101000010111",
      "011011011001010111110011001100111111110101000001011001011000110101101001001",
      "011111111100101110010000100111000010110010101011111001101010011111011111101",
      "110110111011011011100000010000111001100011100001111111110110111111001010011",
      "111100010101001100001101111111110001111010100110111001011001101001000110001",
      "101111110001100100100111001011110110010010011011101110111010101111001110111",
      "010000000111000000111000011011101101101001010101101101111000010101001111010",
      "011110000010010011011001100010110001110001110001011101000001100100010001100",
      "011001110000101110010001110100000010010000010110101111011101110110110111010",
      "110011100000110110000011101101101101010111000001100010011111001101111010011",
      "100000001111101011110110110101011010100001000110110101110110011010001100101",
      "001101111111010010101010101000010100010110010001101001100010010000111000101",
      "001010101111000110100111001101000111011110000001111011101010010110111010001",
      "100010011110010101010100010100111111010001110100101110010010111010110010101",
      "000100010000000100110110011100110000100111011011000011000010110111010000100",
      "110001100001010100110010110001011110011100000110001010111000100111101010101",
      "011011110101110100001000101001010011100101000100110010010011110100001001011",
      "011110110100000110001100100100111110110110000010100101010110000000001100111",
      "000010100110010001100100010101110011010001110010111001001000010101100101111",
      "100000001101000101100101100110101101000011011010001101001100011000000111011",
      "101110010010000011010110001100110000001110010111111101010101011101011000000",
      "000100111000010110110111010011010101001001111011100001011011100011111110001",
      "010000001101000001001110010000110100101100101010111001100100101110101101101",
      "001111001110011010010110001110011000101101011101000110000001010100101101001",
      "111010100110111111100110000101110000011000110010000110011011001011111111100",
      "111011001010000000101110100011000010110111111011100011110000110000110010111",
      "011101101111111011010100011010011100101011110011001111010100000111111101101",
      "010001100001001101111101101000111111101011100011110000011100111001000100101",
      "010001010010101110001000011101100010100011101110111011001000111111011110011",
      "010011101111100110111010000000110110100101110100111000110011001100111110000",
      "101111101000010110001100100000111111100111010001101001000000111101110011101"
    )
  );

-------------------------------------------------------------------------------

  -- constants for State permutation for RMATRIX
  type INT_ARRAY is array(integer range <>) of integer;
  type R_C_ARRAY is array(0 to 3) of integer;
  type R_ARRAY is array(0 to R - 2) of R_C_ARRAY;

  -- number of columns to swap per matrix
  constant R_CC : INT_ARRAY(0 to R - 2) := (
    2,
    1,
    0,
    0,
    4,
    3,
    0,
    0,
    3,
    0
  );

  -- columns to swap per matrix
  constant R_C : R_ARRAY := (
    (
      51, 53, 0, 0
    ),
    (
      52, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      51, 52, 54, 55
    ),
    (
      51, 52, 54, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      0, 0, 0, 0
    ),
    (
      50, 52, 54, 0
    ),
    (
      0, 0, 0, 0
    )
  );

end lowmc_pkg;
