library ieee;
use ieee.std_logic_1164.all;

library work;

package lowmc_pkg is
  constant N : integer := 128;
  constant K : integer := 128;
  constant M : integer := 10;
  constant R : integer := 20;
  constant S : integer := 30;

  type T_NK_MATRIX is array(0 to N - 1) of std_logic_vector(K - 1 downto 0);
  type T_NN_MATRIX is array(0 to N - 1) of std_logic_vector(N - 1 downto 0);
  type T_SK_MATRIX is array(0 to S - 1) of std_logic_vector(K - 1 downto 0);
  type T_SN_MATRIX is array(0 to S - 1) of std_logic_vector(N - 1 downto 0);
  type T_NSS_MATRIX is array(0 to (N - S) - 1) of std_logic_vector(S - 1 downto 0);
  type T_RS_MATRIX is array(0 to R - 1) of std_logic_vector(S - 1 downto 0);

  type T_KMATRIX is array (0 to R - 1) of T_SK_MATRIX;
  type T_ZMATRIX is array (0 to R - 2) of T_SN_MATRIX;
  type T_RMATRIX is array (0 to R - 2) of T_NSS_MATRIX;
  type T_LMATRIX is array(0 to R - 1) of T_NN_MATRIX;

  constant K0 : T_NK_MATRIX := (
      x"fb126337ed0ffbf2e4389aac9149432e",
      x"a216877dc9614af485edaa32f8f9fc28",
      x"67b0aec751ded3c7fed3b03634447822",
      x"1ffe172d815e9eff9449c29f8d9100a3",
      x"124cbc5eb7bb30248d95333a7e9014ab",
      x"ab8df29ec3528a45f515863b4b6cebd8",
      x"67aa2a15203866be7740574fbe22c4d8",
      x"0012c7b7d61b5993bed9d6476a0465a8",
      x"4547ea59e55c31b5686326707301fda5",
      x"1921b4c7fcd32cd2f302693fcb3ab4c9",
      x"13283c51db8b4bb7667db6e8f922a7bc",
      x"940d6cae905019d5153814bfa1f8b488",
      x"cae62c1a9434247e2ab99722ee59c8be",
      x"df7226935c6d09fd1de9e3922b268a58",
      x"6c16fd1887db4f0e11ceaecabaaaf5cb",
      x"c79611ee55a26e6c005815f825d49b3c",
      x"43498ed8f5c297e0502d5a406a1e6c50",
      x"cc583650117553374874594e66db175c",
      x"aa44dcdab477cb6769591483ae9438db",
      x"a44ecf9fe772f5eb663e256d64dc07c7",
      x"91dfc7e9651fdd64f9ba26632bd7dbd5",
      x"2d25b07947adfe4c10845f4650acbcb1",
      x"f908ca1ee240144e99c8ed66fd1b1316",
      x"9a103eca8cc6143c6677b79ed93eefad",
      x"d0226093e30063a930561820af6370c8",
      x"d112abfde53efb6fdc7032ed10c8ce11",
      x"d1caa04dacd7ab1f65e90851e18a3606",
      x"797f81a6308d057450c5d9b1029e425f",
      x"c4174e16e1c3af85c13fe8315df66c71",
      x"dab2eb8443a0e0a169eba6668472019a",
      x"f1a547aefb8b17b5077be24d1fab367f",
      x"7a913da94dc25dd6ae5a1fb1c0382345",
      x"3a3b1e7b0e91f8b1b874ea6fcc0bddf6",
      x"a16f6d344ea82e581c9f5862f65160cf",
      x"9b564bbece1cdb8da0b366a6d36b5c24",
      x"ac92cef46f6359607f138f7d9260372f",
      x"c36935b703ada0f862eea1cb0bd36b7b",
      x"1b3500c999b03dd3f2eccefd9bea35db",
      x"7333599d72ef122b108b52d58288239f",
      x"8848c586c7ee526d885fd16d3ae55954",
      x"77c2cf5adcfcd8e261f2add2aa4674a5",
      x"4b4e746a6cd6b5b0e06c89adfa004203",
      x"d8a73df034c0b2a5ae54a95ab0cfd34e",
      x"7129f8a73213b022fd0d02b470d59a11",
      x"b6aa121739c7e845eadc3db63ed29daf",
      x"fb63b0c719e8e3561874b9bc7d43b785",
      x"e61854153f346f9a13942cef20d2723b",
      x"155bcac97153967f00115048603bf1ae",
      x"877cb6a8e89ca3cddd2a562de758a5dc",
      x"185968989c1d86b25cad3c34a59b5419",
      x"af1dbdb80f5daed18cb1f2da9a99d8c7",
      x"dac33739271995e92180253961730f17",
      x"18a78da5cfe4b173e61c884b6980c77e",
      x"1facfc3609902cfe25bef826fb636b6b",
      x"6a744c36d26f6798ded507b05a770881",
      x"869ecce165d6f507fdc2efc40a9a6df8",
      x"99621ab0a3470976b2eead2b9fd83e81",
      x"4b6451eb6d67b9a3fcef89a225d68563",
      x"148dd7fbdc1ec30a87e037fb0b5f8c0d",
      x"ddf0e8d97acf8052b28129e275324db7",
      x"a12ee70f29635f1ce3857157feb9ddff",
      x"42498baa4706420d03daaab9ddd1716b",
      x"6d5233d6e214c6cd86fe99a70e617e9d",
      x"d80dec33028dc58a1a5b70acc767e8c8",
      x"c49f9ee9258e6d10bc6e371879e33f52",
      x"f17a25f6b784cc1df80e5c5c45adf907",
      x"d7774eeeb2023df7b53e265ce3e7df69",
      x"ab24cde1d3efc82d4f522d7dd904e6bc",
      x"a9ac5f83e320bc129bef20f9834506aa",
      x"d9586b72bd7a6e11e9c1c5c05c35377c",
      x"76113a1e7eb738c6abb4b38f8f35d628",
      x"f1152f66ad2d4d6893b66b89b7f036e7",
      x"c34e163b5df24aa9f77ca933428d6b87",
      x"1f227604ed461186e5349b31010a3a81",
      x"eaf3f81da6390e624975e396809984cd",
      x"0baed6fe121d178e155b6bc5e0530e04",
      x"b094ba94380726a06fe1569cc15037b0",
      x"3272f43bd5a707e262d9a8607d326836",
      x"74c4b0a12413604f70c65911eacd9bea",
      x"e07204bdd0d4a156adea009f6c6c1bf9",
      x"a94e4c665ba16e6477dc3402011d5624",
      x"e2842ac82c32c258993344326950914e",
      x"4e95767b787bd7edac11da37431eeaeb",
      x"875ee0dbaaa5a2c086e02dc09d40bda0",
      x"528f15f12fbc6151782309ab7799d35a",
      x"3fa1b6bd90bd41c2557627ab1a51425b",
      x"9463c9b69af14fb9c8ee7de0df78239c",
      x"1f0948278fb4b545ff87b4ecf3bd4d28",
      x"3cd8722b811524cf218a68447a40046f",
      x"c53d438812d2505713c3e6bf0bedae3f",
      x"5f417dae0d24c42eac7fdf162a3dc30c",
      x"59eb2b0c35894dc8af82412ffc39cae8",
      x"136043192d7b535bc180fbe50179ee3d",
      x"bee3c3c0f8a1929315c4718e5f11a4ad",
      x"e9f65681d1f4df1900da0f0bbd896b5e",
      x"30f583463ac6e1b57fd8c961d82591d9",
      x"48117d039afcbc2f8f8d20384f20bb24",
      x"3ee2494529841deba51f588fe58afeda",
      x"4e24162730965863d383e751489c358b",
      x"a922c1b6abfde633d8b4972364632e7c",
      x"ea4bbb24664639c8f69c2ad82c2942d4",
      x"3a18d07f2583d80ec0a7d9505f059aac",
      x"014d0eae53b7deb42987d554ff9dcc96",
      x"5b022239191054a5f9bf0dd0ea492015",
      x"726f052c760684fc5f8685ecdbc9cd99",
      x"75a77542d236a0a9987a180734610aa4",
      x"6899842c62755634080bc87bdd498a14",
      x"d93abb98c1a05eb027549b6906fef167",
      x"f1b5230ecac6986a02183f931202b470",
      x"a6eef93fcea9abff424faba6f73d2582",
      x"fd0e1037f88c0599a74f7e986bbe21d8",
      x"8c5be1f28d86ebf70c44e62e11b645a9",
      x"244e2834c29c1c87ed012530b302f7af",
      x"c347ae2058341fe84f76b117aa42dc8e",
      x"7363bbc6d29ae3eb58ce76d3f1f1813a",
      x"503ecbc90405f13a84c34620c4081ad8",
      x"4931fb6a84b25f8afb56d1515e3002b6",
      x"4d95b94014e1127a4c011fe406382446",
      x"a8c156ea081feec035d3650fbf454a18",
      x"658715c518fd0cd544d121e1c4f1f38d",
      x"3c2b1683311a804128c22273d9ba3a82",
      x"bc51ce30cab9ab8ebbfba740546efaff",
      x"910fb2b3cdd0ff0746a01e1ac630ae49",
      x"ad771374a75d78344ccd812b1601e0a6",
      x"501bb443ae45feb672f3dc4d68ceaad5",
      x"a3563023f7868463ed42a4feaf6ce75f",
      x"218c997316b9c3c5e6da4ff0f21320d9",
      x"6ba789fdfdb5e524b0b76898156f090e"
  );

  constant KMATRIX : T_KMATRIX := (
    (
      x"d69a7d0500f0be1a0afa96e582f026dd",
      x"ae0a095093afe4ed95996a75b86eb0c9",
      x"0f8531f7e9241696fd6310ea5d69543c",
      x"efa75ed4a280b683fd71c13b6661bf2c",
      x"95e965a594363622d7373e12850aa9ae",
      x"2c5e1b0fa9bd45cde1230e5bd304da0c",
      x"6afb80843997b9084b6dbdceccb1b9b9",
      x"f36aa16e2dea00e2a890e7613822e79f",
      x"32e601749fa50ebec137310dbe514ca5",
      x"778cd8353d2242ee038dd5177b470ee1",
      x"60510da3f88fa88ff6329db8e6aaaf16",
      x"96b90215cd7a170d88a42b53275cb49e",
      x"cb4602e8c09dd59fc2e6dc65bae8c849",
      x"8aa6eb5c0641dbd2fffe61dbaf4cbede",
      x"8ad269a1d26132864bc085b0bbeb1dc7",
      x"fa872700bf4e227e127b8b5eab61445b",
      x"026a0fcd87d925cbe6b229e38753e3e9",
      x"6548e2cd4aada59c6a00ebac06d342d9",
      x"ec96dda9184a22ef9f965f16f6eea039",
      x"397f58124beb92021c91ba96f897c564",
      x"b3336d000aacea0a8d3feb02c443e27e",
      x"03d55db43d653378176f2a9517e3bdc7",
      x"d97636960b197e12ff45eee71eab8cf1",
      x"7f6afa34daa96ee91108b1d613fe0dc8",
      x"bb9b240fe97001c51bcec49263c16b78",
      x"ce736efaea748a0183c04e4698108464",
      x"b22d36df164236731799c2f154d2fe9c",
      x"cb6d5c81ccfecbc62a2277266873b030",
      x"f2c7e8fcb8288c835eb1857fe2150b4f",
      x"772a7f35934d569ef4b44f271e420bc8"
    ),
    (
      x"683f6478b263b6df257f67a44eebe296",
      x"168e2195c8ac90c203c95ebbd7b92803",
      x"5ddf08bfeb8511cd5807057c5b19078c",
      x"648fabed53712496e63295e39b060d23",
      x"2186d2ff74daea46d7c2b84d47bd732d",
      x"467727e023e7babf087f2cd7364dd4cd",
      x"7f4ec44132a6da97dcc28d9d71794c5f",
      x"b3818daae8a76a522b8cee68b3df5c16",
      x"585b5d2fd7e4d3079834a2ab9d0f2a48",
      x"a3a06ec87da0774095ddefc06d72182d",
      x"de6eee1dc27156d0be95becc913e346d",
      x"00028ddb25d316c29017983fb4925410",
      x"5c2f4b9ff9749b7e445395e36768f6b0",
      x"bf3936e7f70b903fea635745109f6e5e",
      x"c2ef460f65d8edb1a46cb24ed89f65ee",
      x"d4d0b779ff441a9e272293e3f241baf4",
      x"c8b70969ae36a41ac8d4bb23194d893d",
      x"e8ad0d6fcc365d83db9338a60ca1f592",
      x"23f20ab7f70ae73c94d39c57dc3b332a",
      x"863e4c41be196d47be9818dfe0f62f91",
      x"fe71b032e634146bde3d8f63f2dbedf9",
      x"893b07159416c400f60f8e6faabbd2a6",
      x"646d363743e559b96b2f7043ea197aa3",
      x"f1c92bcd47cef88957cd370ecca15ddf",
      x"18d5866571c46bf32f7e8d4bbfd95365",
      x"34d13f9441af09b7dfcdaef45f7a8efe",
      x"a6aabf25e8854d060a9acc3a69d0fe70",
      x"50262be21f9fcf0c0453e988f30fa00e",
      x"125c9d7cf069060fbae019204e5a1e14",
      x"a43702fbe370963ef36c75d8a8b6cf2a"
    ),
    (
      x"676633d87c8c6781c10bc25ae6f75878",
      x"5961adb11b7d30ee7b499fbb41b7b4e2",
      x"47c338e1beb9d93482d31165cac78547",
      x"cae832b4d2388495a528fa2901cf47f5",
      x"40913daf1d44bc32d04fc0e6241a0d18",
      x"8e1aaad8dcfab9029249a362e0c3afc0",
      x"7e1b96b1bce08be5d4efc5944ed90ba3",
      x"fd13db9add8496b80c8e638f8d4f06e0",
      x"7ea9f66a4364d87c82aab648d0c8e2ba",
      x"4a9afaad839c4a8090cdaa9febdbb639",
      x"7a8c0d2dc3dd4a9d6dd7d1074004344f",
      x"3fb9bdb9ef52c1ba91153e3e5800bbd5",
      x"b966f449ecfafdedb5e2c2b71c379d4c",
      x"da4d6c1ff47740838b4ba600d8ecbed4",
      x"4e78424f70bb720243feb33e7d4c59ac",
      x"eeb24eb6343a0410b832eb620b3dd2fa",
      x"011532ee86336424642ee378e4fdf774",
      x"2adb2af983da0ff53c2e3f7b8a5b22ce",
      x"4ea8bb5c8bf2d397f44cf95ea0f480d7",
      x"4adf8dd9eb1ad7032b05f9915fe8dc11",
      x"606fe2b6ed3a07eb5f362583e9e71ed9",
      x"eadaed902f07b1dc74439183dd3171f6",
      x"35960075bbe87f3d521651da1146880a",
      x"09a6db7547749ec9de5b221e6ceefa72",
      x"d086c33a539a369fbf087e4da5ec73a8",
      x"71746feaeeebb86f797647ebb947a40a",
      x"6e0ce5d8493c49ff213407b32b81692c",
      x"98974bf6aeb99a0cef6e0db4da4adcf6",
      x"8bc507139b7e2b8b1cb484e61c7cfaa1",
      x"9af75b7e1a9fb3de1a4d4352ccf30449"
    ),
    (
      x"85ffe3eec111c19d8a8f7577d17ce43d",
      x"66e6cfba729a12846fb186ba7da1942a",
      x"6b01282ae106097a7e090f7cf0672698",
      x"06984683c10975970d70ead0e1bc6f8f",
      x"bfced29f488f8b6b448a1e7006c2691e",
      x"8afce995bd7863829c1152c982f35e3d",
      x"6e2de74db0a626c5aaf91a76c512086f",
      x"c3f953049cac9c0fe32805dd9776dabe",
      x"bbab7b68998e4f02b2fe33f56f2a81e7",
      x"1841daacd7acfd1720d1b5fd36f0c18d",
      x"1a63c8a88c3e326e2e1de0520f9159fa",
      x"cc84e6d994e8b634a7f9d8b4ec0e9a01",
      x"d262ad074530b1284c68e99a913454f8",
      x"5c289b25059af1a79839e90cef4eb7a4",
      x"dbb4c22b380a05e8d800953fe41909ea",
      x"cea3f3bb9e79b03b491374d6b207a15c",
      x"f3f2f20ac8328ea1bdaae36ccb060d02",
      x"492fba54ed1675769b063c17802d36cc",
      x"94557cb30b4886d38ccccaebbebc7b78",
      x"a98bb62cadf4abc40b8123ede9382459",
      x"7769005101ee7df0fb6decf425d74cde",
      x"7f6cd22bb861526abe6dbad97d42cf73",
      x"878c0e05e0a6861d52a095fe1b1260fc",
      x"cc05a0290f48e38afc285b0bd49b6082",
      x"b086ce239af16b1c993a71a872a4417d",
      x"ddeb7edb5059177136d3c26be63d39c3",
      x"3c7ca7b05abb1444672a8dfd7fab05cb",
      x"dedafc271a9e2574590d388edfb5ab94",
      x"d6b924a0fbcc4fa8a3a3014b25adc5c9",
      x"83d1d027d4c4908ec53ac8eb132cc8bb"
    ),
    (
      x"449ce29accc0eb8bf13d17deafefa5a4",
      x"99e888e308903ee8bd13f0f4d8f026b2",
      x"0e29cb2fe7ec6fa9529a23ebc6cd8831",
      x"3c5957c28db246e62e1758f93e9d549e",
      x"e845863834f668a55bbaaa101d21db3f",
      x"c8278b3b3aa22640c6291ef5fe387080",
      x"34e896e0dbf1a6a34acc2781968354a5",
      x"a7e27de05a0a532ddde2b5736705ac4c",
      x"ccb56ff2d2ca3219b2614b1e82597110",
      x"14a50070b9213830ff3377fb893b4bee",
      x"ce1f0b58a60eccf549f283d223cb319a",
      x"b10efd992fc51878c3b8e2adb6e73ad5",
      x"3e99b351469731df2a105026a6fac996",
      x"5227bcc5f433ba93e2c5aeef63f3a592",
      x"4396817c6f0fa9a3668d0ecbf5fdb775",
      x"9d0a4d4fabeafaa10f923065ff654c70",
      x"53a48b9c65200320d49e18366ef66cbf",
      x"3d35d5db79f98287285aa0af62e84ae9",
      x"55c585b2c7a2a5b6a4e6f3930a059843",
      x"4fbf4ac2865e533d9146f8e9d51d216a",
      x"55486de363c79cbd74c42201115d4bf2",
      x"94940ec1b821ee1857f9293548ed015c",
      x"a08cb63c02fd54387cba04ba63b1c372",
      x"28c6bad1b70802b5423abd8352bad8c0",
      x"2aafb420d62b3c702685734ad12bcd60",
      x"1b002a38f85fadc93be1d8d9226f99fe",
      x"847b57ceac965db4e559cb0e796c03e2",
      x"eb0b2a499f0f98383317b4c7dc616cef",
      x"4668fd1d6844fa9037cbbf5dcdaa1e7d",
      x"54a73d0ffc109e1c03841a7b55738223"
    ),
    (
      x"0d47faf7b2af1211ae4584a1b2d2a91f",
      x"98788e38a72eca1c4e37237235e99c89",
      x"a8c9e5809a397ace898de4d285ac0637",
      x"75defb7a31e1896fa78573cf783b76e0",
      x"6a1e740a8472403f356c94fb0f41c794",
      x"5bd573aa1949817778e01076bc8a2028",
      x"8e979149fe363209caf37e2fa3fd9624",
      x"aba32fe9e798551cddb3c7170191c649",
      x"2d93d956e2250c2006431c6af843ef72",
      x"5c3fcd7ef6fa8851ded39339e966a6d0",
      x"ab91b30ba805716936fa62e4879aaae2",
      x"bbbf436d2e7c1e4080399f939e61f5bd",
      x"8d32fd7641f3db00beeb29cccacef18c",
      x"37ef9b42970437369daceca751f10be3",
      x"164ad08a02ac78096e96b74a2f55dd29",
      x"244129305e7974a1401fd8b6a87bfd8a",
      x"97c09f5128dc6b04f410f5b467f3a3f1",
      x"2c6d256dab04ece3ea96fb79d598ff81",
      x"00480be984b753451e2683ab4780500d",
      x"58868a38670ff47fd01cc8440a0d246e",
      x"a57ec1bccc2ca906e15ccbba8866a51d",
      x"917ed8c9f7ea81cb410b75ac3d99bdd3",
      x"ed3f6cf73d257ca2fae9421bdff76d9f",
      x"774fb680a06f212ca0c27f1c32111002",
      x"4332c28d533cc394e07cb3226b4b7a7f",
      x"e0ef58acce720db2551bc82791dc9487",
      x"6e8da7c7ae993aede359c9c7d7fa7236",
      x"1a9384fc027d2d38a08b3a44e3d957c9",
      x"b65f58573705711266789d9aec296846",
      x"cebf85a3a9b275fc807aebc0ad5cd845"
    ),
    (
      x"128e9f75e67563bf05cffd1503d8680b",
      x"01deea243bfde1933342b3b905c50e0d",
      x"ae22187fdd9fbcc2826e3da4fea18648",
      x"23b19d43364ba21b855934b0ad9cd677",
      x"00dc46e0f78706c514772e48593ee170",
      x"7ebad13f93555203818d9e0c0c9e2f29",
      x"6149454b4d317f3d368b2e8f18113686",
      x"dbacc37e44d9116af9bc0aa95f72e0f9",
      x"e9df559c426faaf943068368b61cc1ff",
      x"a49fcb21a3285473d94f4574d3762f71",
      x"90df0ae68ade01368048ed6b6099f380",
      x"f94f93e7bc214c580086efca1032a373",
      x"7438863db3eb4a8a059d1a02da6d7a52",
      x"d1ea25e580b8e721c2d64c58a1188067",
      x"f14663e6bbaefdd609a790e0c20a06f7",
      x"41a10d8a0134e51ffb7d214eadb194a8",
      x"ac177475bf86051dd2643dcb87c49ffc",
      x"9527c3d03877b3e52f9eb3d18f256f9b",
      x"6b454f03e068478fe3e3147813353160",
      x"c280dcca219ffeee538f47a2f307ba63",
      x"01b99f897421a8ebacf7319a438a9d75",
      x"748a93c7ee6605098ebea3aa00d7ff8a",
      x"7edfe9a9b43370d02a626885a4abe407",
      x"2a003dd8141ff6e2b4a94b259ae92141",
      x"1a8169dda632aff2db76c429d0e4047e",
      x"559ea5b6e8145aa865f8fcbdc2d17dad",
      x"5276951bcae5a2bc77bdab11926de924",
      x"cd20993cbb7e8393593a08d2e3b18a7b",
      x"8a74f20c78f64ef44809f6a2a19e110e",
      x"42270a584a9d92f6ca0798e5300537b9"
    ),
    (
      x"030e0e8c5d01d887df1e3885e368a2c4",
      x"51adc6cb7b5d561650dbf58ceddcae16",
      x"0d7eced06682ac652f77b8c235257e13",
      x"4dfa3e6701bedb30a24209605b15e67e",
      x"9ad525dfb762d4074938a703432064ed",
      x"de1e4050f2e81a44f2a5d2cbb95536b9",
      x"ee79dc25d261c5aec1810ef9055ece57",
      x"9b74e2daef8428e968a72f781766dab3",
      x"a4ef2ef91b1b7940452ec3cf2470bbfd",
      x"a13870210526041a3a6478ad9365e35c",
      x"b08b878a2b6497a0c93bba3d0d44ea22",
      x"d567077fca7e7ab4ac367e900b8cb4d0",
      x"b223471f1f7f2c84a4753bcc34cf595f",
      x"8464e8369db8b290740bc5fa2ced05bb",
      x"e4cf3f741310d71c1e3bfdd36fb4e9e5",
      x"ccd1520fcf3b1619612b20d1bd57fa2b",
      x"51b19285ab8da25bc438a4a96ee97fbe",
      x"c06b0d57d8b7fd0aa5d598f68e146233",
      x"5e7670a7759c5940b9870f3566317fcd",
      x"a22db34d974c3297ac197b42529709a7",
      x"a4da2525327a0618a4a1b5b6b863dec8",
      x"021b5e631c6de7f89dae3792de842f2e",
      x"b7b3b6bc827e8d6e891e5f47d63464b4",
      x"3adc5eeaba21a35901a8b57f0c96cc5b",
      x"36f37c97490bcb3d27cf12c44f23ae6b",
      x"752d00bafccdd9490e8082aa5c818607",
      x"9758ab867851e2808e2d3fda80c17cba",
      x"d72a517ce79f2a0eca7e3c03ccb3d10c",
      x"f3f7334c0f525d9d8ea1d2e1d47f6b54",
      x"a912fd79c578bfaf886813e527c861bd"
    ),
    (
      x"26487ce0601d87e879df70f872745983",
      x"2b7cc61a172b909f2fb60e2eb312c42a",
      x"078c438e1b7ced0c058554f77d7ac9f0",
      x"2eb2063adfb98cb6a78e965eb7a9436e",
      x"ba30f90f4457f84a73767de55a188779",
      x"0e029c7b8b62d8fea3febe0ef3ac1877",
      x"a67a5e120213743303e584e55d6991ea",
      x"e944f09ab34d4ff6338272d7f487b368",
      x"e0155e0480fc78982f6a301e6b8da3b2",
      x"5d0d648ef30a381c5dae8c7e0bf13935",
      x"8f235d72af062ef57cb2d9477fe8825e",
      x"438604cefeaabcbc6529de486b44d0a2",
      x"eadf3bbb85ece44c94e57b412b982e15",
      x"26d61367014d044f6fd1e7ed9126a19e",
      x"ab8098a2fa23fe5116352ce7354f48f0",
      x"902281b67390b7c4c2042cbc2c2ee165",
      x"95c309f0bb16c18a01c3d0e50f525080",
      x"d276042ffe7af1726bce1325975fbc3f",
      x"168819c1cb7d2bf3260964bcf5892e03",
      x"c88478fd88cf9ce8b69462a8a4052b38",
      x"7950b7ec1a52270d9ffca00728343e47",
      x"43aedd5391d0a5674812a7d400f62871",
      x"348cd20f256515f33c9b06aac253605d",
      x"ca12c00512c91f4717d734ed852dd7fe",
      x"5279a1adaf93f8be1dcd3bbdf60782bd",
      x"6b329dc647f664bdf9eee11e9516795b",
      x"e8a12f9a7577b77c1cbcb4c40b1cc9bf",
      x"2941b4a9e8379ccb68ebb032bb7266ed",
      x"9b68f868751338ec0358e99764febabd",
      x"da9a807ef33e6b76abf079027f508695"
    ),
    (
      x"4a7f57ba225d641cc91f708b72df7e0b",
      x"b17a2f9591db9caf6d6d75f8825c935c",
      x"01931fd97ca3791b3dd2bbbacb62b150",
      x"fb442e9b482fbaecec26e42d622ef8ac",
      x"048ee142191e2d2b75cc5df4f49668c1",
      x"20583a036d1887d0c3e798fccea05f02",
      x"ea4284f911ba01178a8bc5964a608b87",
      x"150749abb616e28f3161c9cbb0c8b3ae",
      x"2c0978b1e8f77dc5e02eb740c0f51bf3",
      x"81ad9ad1c51f0bdf0f062db55b8f5926",
      x"70b7b707423d777558c59b514054462e",
      x"db124378730b04946ce94d3533fb9fbd",
      x"47f9bd6476e0901128304294dc6a6825",
      x"e00b57603a6276a5c6277789089675ea",
      x"4c318f138d79e40ced3990389ddf485c",
      x"571c1487d87166f6faa3544cdd8b086d",
      x"70c989815a3d23d0a6dd9eb60c2d48f3",
      x"f5a59d02611e350c28436a04ee00389b",
      x"a9a0e4c88abc80c12e4a1f7140536cbc",
      x"6ea79ba7ac2e17d02374285c0a3a8582",
      x"e23033749464d60449b9f98bb0ee4565",
      x"a9d79b51ff39993a3ca4f5ff99bbe0e4",
      x"d8a3ba459c7a8aad2bfaeb275da29757",
      x"532b3f3093ea93fdabddb0212e2f18e0",
      x"80f5e40870d9c4a2c4debeba2109f8cd",
      x"be8488bfb46b5d7b51257eff7c2b0de6",
      x"7eb8161640ebea73dd276fd51113fa3a",
      x"2ec5fc7e497e830df0f11aa83c671377",
      x"20deac4a6f20de29a29b438b0940f440",
      x"1c31e52e908ca3af9873592e7e713123"
    ),
    (
      x"5e7541e9aea84b411038e8c941d415c2",
      x"4b355124d22536866b2539766db68c12",
      x"4ef71a79f4e1e60f90aed39d51af5d43",
      x"7ee98ea072687dfa1485205906ef7ea8",
      x"743afe57779b276be8058a867d49aaaf",
      x"a4660096425d5b7ebeb648741e471bb8",
      x"95f32e30848bb9fb5ee93a83f597db33",
      x"58d4d61482dc80aa7203d2eecdc7aac7",
      x"2167923c8d8541caa032ec0493de97af",
      x"5723d5178c072f87bae72fc898f4b0dc",
      x"d94d3620786ec17254ca650e816066f2",
      x"33ce113aeb35606a4bb6064a9b352b45",
      x"f3a0d1f41cc6393a807e59e99bf15758",
      x"b3bffbfb9b90529dd339f91937d93517",
      x"6242f6ad0c18173be80324f6ed0f8f92",
      x"26ceacc1bd5643b70a81e1a4bb141a18",
      x"80eb232e43de5f4722f3a2f05a74575d",
      x"e29420e773707483414eeacc0ae9b6dd",
      x"2ecf96b1aac8288776105ec5699c200f",
      x"767526c1c029ada057c6a3a0855edac5",
      x"bc4be4f6cdd1f77bf6494f8bf5246542",
      x"db22e0ae80fe29cf5ec50a6591242f63",
      x"cf1df75e32f760b3138686855ea83103",
      x"0aaa673fbbfca4ccecebc8c9c77e67fb",
      x"9aec755db7aed424d4c5876789b7dabd",
      x"5c86a00fbc4883691fc5fd8ab6714f76",
      x"45e028b77286095f347659f0c33f5f9a",
      x"ee803801dc40fdb33bef6bb45aa93146",
      x"42e0268c41ca18f5ea07ff3015051285",
      x"6e7ab42108015712c23a314b63c4c2f8"
    ),
    (
      x"b59c2fbfe36be28fcab0e989cfe84315",
      x"d060647636a0ff9400a70ca3436a852a",
      x"b445fda3d4a2ae790da9a30d6844ec15",
      x"03a73ea5b2c4539205c326d3583d3e9b",
      x"4ae7259cdc6af65db1d1ff1765805098",
      x"71970f21ff28622564ad79820ae62ad1",
      x"8c6937bc82dfeac6f6e4ee55fb73e5a4",
      x"3fd9cf593116549e045514e41c004aa8",
      x"605c9342e69fed2baf390f3006671bf9",
      x"5d74697451b414d7f27f33adb8078300",
      x"172aba03abff8b07c4e9982ff696a821",
      x"cedb12025f4bfe03ec597240d469ff98",
      x"26a1aa6c4a02c1baf35bdaefb50d7dce",
      x"00bfd974e8e1497f6934cb46c80fc693",
      x"09b568c770b49781be1383570330ec26",
      x"0de7bc3dac27fffa171ecefca24effa0",
      x"39eb1a2e122fdf3a3f167d112d7b8fcc",
      x"9c85b9c3861d2850bdd2c88ee4286b53",
      x"14df7309389ec311f3825f0c8b5e5b08",
      x"f39e8232dcd94ff5c284106667fc3106",
      x"721cf62bc47e2b3cd5f075848df89248",
      x"6e48327fdf7c372b7b737f832210e3d9",
      x"97557d07cd0e74800cd1d379f0f8d05f",
      x"7d261f421371a375d5f28930510cd4d8",
      x"35aeb085d9470de9d72d7d640ac99a5a",
      x"bffb8f674a96bbe8c61b5c09249dcee6",
      x"115fa96ea4ca4809ce6fa86e78268241",
      x"d5b84e7fe738edc81d1eb1614b945b7e",
      x"1d6698603b50562c35cbf12dff2b91ef",
      x"80b2968910889aa0489e7dbee7d01d8e"
    ),
    (
      x"bec1540d39a9c80c1e7fcd1a7310b39d",
      x"9fa383df3e4bc61b1bc24f6e32cea283",
      x"563350313e7e6753c7aa79b916bbf8f0",
      x"2c7e6136b2fc1aef53407f15295dfbf1",
      x"be9a67a809421884a9ddad24fe494f64",
      x"f8bf39c32522ce508c9175ce2cf2e269",
      x"b0b12514c04d082703fa1b7e2932bf78",
      x"600c49968dc3894585508076613ecaab",
      x"3a703a496a4190dd5c50ab645afaa80a",
      x"174155a5cabc7d8a270e0e87639b7d9b",
      x"a5fd1cef69af0f2a17edc47f5900dad6",
      x"3ef01ccdd474281e4a9332d4b4bdab80",
      x"78f836a628dba5cd272cec4432fe9309",
      x"50eb2f21f18671676fba623fd51f4f1b",
      x"2e31b3528be10f809afd3c58fe0ca4fa",
      x"e059dd23d48b60b28a4e7a9ec30806c0",
      x"44ca9da75aa76d85b3872327770ac54c",
      x"ffcae2c51c8b01e95315b1ea51bfbfdd",
      x"c4443b2a53d1befc25d6e8dec60a5c3d",
      x"2c69f869fa8c63b35a0b0b8a567426b4",
      x"5feaf433819b8e998ce3dc8416558054",
      x"6d3af8aa558e2e3155139769bf76bf9a",
      x"33a1eb81b41aa5fd699a6fdded655116",
      x"1e3ede616859792803e9f018882e9aeb",
      x"7570123a389c46c7db3e67d6bc684d39",
      x"f3e0585461af168aace299ed84cb0a1d",
      x"766d3f86f01ff0b9372b30a8ce1d17ca",
      x"232455e5af116aaa83d6aada3c751ff6",
      x"5ad0f942af87ca9c5184c73a7ba58729",
      x"ab6878aa946f5d3ca772ce6ea2d00994"
    ),
    (
      x"83f432ef1d3593287c73d18973c733b5",
      x"1b7e10067cf68ac0ff4c1abb3c202ef5",
      x"d431d32356141ad0a24d9e1958a2c816",
      x"de43624b6bf9326a47ffc656d0409ecb",
      x"d922024d66d53190198d5290efd6bf75",
      x"066d7b099186d74643cf8de5eebcfda7",
      x"3950da988336bcaa50fb10137a1a9407",
      x"1e7a4576f7a8bc2d25f6547383aeab33",
      x"cc7a46f49b0ec8b1a8c3b32257f742c2",
      x"0e0632c89796177ba33d1c14223b824e",
      x"98a35d0f1688f006435e225998b01a2f",
      x"e04ac3bef76d672590f1ee494193c4f4",
      x"6f78b8acf703dfc3ca93c04cfab7f119",
      x"9831ab3952fc42bb5bf8b08fc9d7d14a",
      x"f5de75a58920832f8709d03627a8a722",
      x"52455f3d22f4f2a471ef9c8e4ce10d4a",
      x"69055ad9a0c57ee22f3e39307b5a48a2",
      x"7bc913819c6c20871679b33471df7005",
      x"320a5b2a23e2848e00502cd6737a559e",
      x"d5660043f3ecaf1bfa6003b5f2f75033",
      x"27891bbaa1d970b9a36c969fc35e1de3",
      x"5790aa75a0034cf418d686e7054502fa",
      x"baaad026113d575921114b8c54b77f28",
      x"219b403f4b4cc26838506a2bd6b5e91b",
      x"81bacaa30b7df93cd9fb9b70c3131019",
      x"38ae1a11fb2d615807bbceabe9d59c1c",
      x"bcc6f3dc9ed54c3b12c3ce3f9c6999d8",
      x"c8ea41e46e7a0c6822daa976feec21a1",
      x"a7e694a0f04b84059ad4ce657af02a7d",
      x"e0db4dc12df6f864d083983c03e41fe0"
    ),
    (
      x"954bafb8292601de797f53517e3a450e",
      x"823ed3dbf29c64d420ce4b9e3df0fe15",
      x"38bf5a299ece2bde222a884d0206e0e4",
      x"ca8215d65dfc082ed9924c863b459a17",
      x"c2e1cab648539fe19452173c0394f9cb",
      x"c6e38a87178b357e4242d308c500f582",
      x"b0fe92382facd84b30245e762c52b6b2",
      x"0dcef2a0dfd4c014c98ae60b7a9d7d5b",
      x"e294158327ca21d6fc10679040dde44b",
      x"b2ac5db5183a9a9fc7b5499db9f97a27",
      x"b2764d70047157f5eef4e6548141e2c2",
      x"bb487eebd2ccce79983474bc74064bae",
      x"460d02a2be3863b35d12eb8fbd513567",
      x"54c3427deba5bfc0f067395b67760f95",
      x"fae961af0eab18c77a60d53d931bc5c8",
      x"9e3461fa86bdbcbecbfa72273c9ced09",
      x"ee266754998db7fb8804b2ae9fa13d18",
      x"be7eaad6b25cf97f758004e76fddc68b",
      x"3123660579582397c2a16f928433a636",
      x"f7950802a1dc4539c9c66a44d03c69e1",
      x"c1aea156d1f21b2aea5e25a391526073",
      x"90939d728f4c9d0e92a35f1cb28f51de",
      x"bf63cf616ebab4006080b82e38a01c56",
      x"e5169db7b0cab99c81a5ecdbf796220c",
      x"ba8bbc1c49d64585d721728acd2231b3",
      x"e4ddaf1b7aa5fad1762cba11a6d32f9c",
      x"bfea3d61f580a16a4b5dd2c75d8f4b4b",
      x"e11013d2794c7f750fe3b7ea2b5286a7",
      x"59adea0a3a653dbf8691b253c602ecaf",
      x"06316d436a54cf82d3eec1f15d544421"
    ),
    (
      x"6deb1a3c6045ffb01c2e1dd8ec8d0fe2",
      x"1f0fe236625fb12712463822b2629610",
      x"87e63a7ed481460e5b98b405442d9707",
      x"4abe6f2d34cde592f23a2819b583a033",
      x"5cd1d3e5e5d1902de5b00d9ff9541b48",
      x"0d8de3edba335707ff65154d7008ed3c",
      x"c1542b357e3b3d5602c38078862025c9",
      x"585380acfa0e378b4e6884671feb0d1e",
      x"6f2f0c720a4ad62a36d7d31f601e29e4",
      x"263da3f58f0a85147d588b49191fb837",
      x"be82eb31f608befdffe3411962d30d34",
      x"254f6f9c9f7d830fb0701cd6c70001b7",
      x"46704d7c1c1f1a759491758bb27341c1",
      x"3ef4b134c57e23fd1d7fb0e61a4da01f",
      x"4e371a6f96de0b29e270c529f8fb969f",
      x"e2b85b03ca15171e0392514693c6382a",
      x"1a085cc6255a1b6a2dcd9e3b0b87dba4",
      x"36facceb38a5a906711e333198da5091",
      x"613147e1add31b2dcae45881da3e134a",
      x"43d3ae11a79d69a42b808b705ee46e67",
      x"724ec048942cbdadef6358c0f81e7015",
      x"1bf63e6503bb30c3dd4b5de0950be08a",
      x"2eb1549080ce1647c1546b5575a334aa",
      x"d892fe95d1c68401c888bb423de10317",
      x"0176a6d8166386cf50c97151ae69a406",
      x"75776f9e4192fa204702256ac4a73b71",
      x"74b20fd3cb52af64b5bdeb5a2c8ac130",
      x"2e625c1f88ea8634a4f1b4fda6def461",
      x"7306dabf2df3cd5e417a5f72f02e9331",
      x"90de0ae2c967a2ef0068a8c7425394cf"
    ),
    (
      x"d8ccfeb0068102f477d0622467208b7e",
      x"5b4538be311e2bb37f3e7cedbe4bb61f",
      x"323634aba39ee77e17a2efced7f3f31c",
      x"556c605daf51b792f8761e8962f6345f",
      x"4ef0e9993f60cc75544f7a16abf70e57",
      x"8cacefd2d34c34a88390fd049a02319b",
      x"f40ca5b93250da86633d8d528dbb8a78",
      x"a07066528676fa246c3f6d2a73f11a27",
      x"d6f7a19cefe60001181fe75de2f02ed5",
      x"b412de6f0872696b33e8110ce8bbe423",
      x"3b4cc927b50a66da66660d7ea0195031",
      x"3817e62cda9a0fab59b37f8688b6b011",
      x"7bcabed77728e78e662c8002b3fbb867",
      x"dd4d78538f15d17c3e63aba56c2b9601",
      x"646d0ea70e2aec8421130d6fcbb31e68",
      x"5a9f19ff933f0d8a722d76036affec7d",
      x"37fcd297d411cf84dd356cc1849c235b",
      x"5c64999cea55f1f8d6dd98cf0e7176bd",
      x"10792f34cd1f968dceb0da2f8202a141",
      x"824a5cccf865ea7ac9c9160171696c3b",
      x"dac3b3afa204c32568d5853f112c1c55",
      x"ccbe818cf0f555475c56436e38c0b0c4",
      x"27a77047bcb7b5e9958195977433a56a",
      x"d6e24dd4cc39705bd7a7c6e16a5ed97a",
      x"a2f0d58d479eb3c032dbc9738e69cc12",
      x"4b352516af0a2fef9025b458537df846",
      x"247c79a48f9c447726b1dae46aa4ec80",
      x"26e89d053357364f665b9dcf037519f1",
      x"fe5ff822b9a9f6ee72119a2c930bfbd6",
      x"73423df0824991a3571aa6ae42385eab"
    ),
    (
      x"6e71275c3920c5237a6d4a2ab5dbe92e",
      x"732e78a0f4296e9bb3eea2f44ab6fdf0",
      x"066df291982e1fc0e5554c4ced0686da",
      x"2365e1f227e7b4af0e566726cce047b7",
      x"ea888667aca04d9064db997c23c8df3d",
      x"e90c3b58671e8d58ef38fafaebebdac8",
      x"a41aba2831dd14029c23591489ed8c4a",
      x"23abfbbb1ee87f7fae3694d85acd5b29",
      x"91f5dc37795934c59a36861d7a0e08c5",
      x"679c6011cb5e66bd4b6d0a25ac8a65c5",
      x"1acd97fa5b05343ae3bd6df95919e857",
      x"2cb1b66f4f87af656be708081bd37804",
      x"0a0ef95a6c040a09813042fb69d1356e",
      x"8c1d14a35aa823aeba93416419039c12",
      x"065193d1130273d07aa29f5c398748a5",
      x"d88e71a20055ee861eecb5f5e316f270",
      x"93438ab61749010b8d35a1b0962fad50",
      x"a5ed560524b23db74f2291610b5c111c",
      x"7db89a5aeeda13c90cf5760be506023e",
      x"205bfa1760ffce282e7fd1ee528052be",
      x"f5928dae61df732a26a69014597930d8",
      x"ea1890a701b31dfaab23763d0bd987a0",
      x"871c6ebc151184e9c7a59ffa3f461de0",
      x"cf69f6dca1d1aed0e3f4002c1851ea9f",
      x"b2214dd8740cc4dacb8107596cf9041d",
      x"e22f92bd4e84a6e2bed3c084c4e6444e",
      x"83c498c905c3c6732ba8a5e8af8d9c33",
      x"b447f9383cbc2491919cd5f3a05d2dba",
      x"511d44535a1469e20d010cb226ac908f",
      x"6e875316331ef5bc80ddc0817632c7fb"
    ),
    (
      x"f5ab0ebb7bb8118d349f5732ec57f5d6",
      x"bfb4d2482e2ac38f22e7f0ce894b0d93",
      x"fb460334d675d210e2fe16b55f284522",
      x"e08077cd2403138af9dfb1647b90e3ed",
      x"2bb4e2061a477e54dd630b014cce23cf",
      x"10e36f12cce8f189d894c1f36f6c11fc",
      x"6204c6a8454b35812d18ee04cddff292",
      x"2cd6b38b97e5a65751943339d6b0c4da",
      x"8f89cef5d6b06d3fe440fdedc217e23e",
      x"0786b34d75a9ea6b89934337f69bb119",
      x"b15600b44bf364369cb1cb54764452b8",
      x"f89ca2bca384ef3fc530bdbb3e01b4ff",
      x"5a83878197ead0f42f6b7f52ed38d460",
      x"d035a4ef987c2e60e0a85c6ea6f6f217",
      x"26b738dbf608833df52a529791d8bd09",
      x"a2d79741ad667174f1ea91ef9c5329b2",
      x"0c8b2c96a3bc61cd7b88d8bc4d13feb4",
      x"0a68eabda6b52707723641bcaba36425",
      x"4fb0e95bc605633533d6c421561a1468",
      x"25f20dd61b6d6c692d0afd5b7e5108ef",
      x"91b925f053654a09a6e2edbc2a7a358a",
      x"1df628162dc27f7d1637549ccd148c36",
      x"754daf1c4969236beb44d595f6f88d59",
      x"d1927054facdc89008f9f0c27f2aafc9",
      x"742e6e2d8d0f66003ce250f8671eed74",
      x"c36271c2d3cff234408b7fd6e457ad87",
      x"35da472f2081a41a8c8c6240de5bc2df",
      x"821dcf20d0f375b2e562999e7a341466",
      x"d821f67f9cb271e1de1555afa8254afa",
      x"95cb93cd5a0ee3413942383f4edbd855"
    ),
    (
      x"d16c343c9f141a870021de9149a03475",
      x"3f6b0e938582dc9f3bf528b0c7213e6a",
      x"526cb22992ec1cc67124a329d12ada76",
      x"e7d65a29ef9974409c6dba3ed5837745",
      x"a90ce717ab7e6c419037232a5817663c",
      x"ad9775af28daa9059be4d66161be05fe",
      x"d45bc3cfa9ed6e8e0066341873266a90",
      x"84afabf6462cdecbaa34aa9dbdd7e1d8",
      x"c64d695980aceca22a2f81a459a45bf7",
      x"d21579da38bd51e7819a68df6fd72df0",
      x"8e8ad6e9cb72e8c7042baa038843d1f2",
      x"040897015b6abd01fb68456ea191a7ae",
      x"f2b41fb5c1906623bc08e26cd0e913ee",
      x"da3ce3aba51c9142cbd0ff30263b6c8c",
      x"0f272cd2104043c9bd9a6b7bab839b45",
      x"4506061266cef9adadd9dfb89d92331c",
      x"60e78e5042b7f9fcb552280ce3c61e5f",
      x"251f53e57d416a0cf86633ffbd890e82",
      x"aaf34b97fb9a98ec948956d0b7990c54",
      x"d13b8fa06f1d1f4a97fec912d1d80602",
      x"49366518e411fdeaa9808041ec083261",
      x"d7ecb020d9cd9d5d8e3db66941877d6d",
      x"e4a941dfc10d8886e50506d503332939",
      x"75a343449555c3f58ecf43fe2869046b",
      x"d3a95bd293628d8de01e595e417e5f58",
      x"48790bfb7c534fc02ce865de89c9cb58",
      x"59ed2e74b64a5419de209acd0fc0b386",
      x"f22dda92be29faed5b9528d2c38fc851",
      x"9c169c9450579868ae5d077e1bb156d1",
      x"16e8de5576ec038ea97166b4385c9147"
    )
  );

  constant C0 : std_logic_vector(N - 1 downto 0) := (
      x"000000016ee016559278ab60a47f1a8e"
  );

  constant CONSTANTS : T_RS_MATRIX := (
      "000011000001111010101010111011",
      "111100100000001000101100000111",
      "100000001111011001110111001011",
      "010010001011001000001100001111",
      "000101000011101101111110010101",
      "111110001100110111000001100101",
      "010011010111100111101001111010",
      "010011100111101010001110100000",
      "111101101001110110111110101101",
      "011000001110110011010100010000",
      "011111100110110001000010000110",
      "001011100111100101011001010011",
      "100110100010000100101010000001",
      "111110010001100111101110000001",
      "000000011011101011000000001101",
      "110111101100101110011011011100",
      "010111110000110011000010111010",
      "110010000011001101001010010100",
      "101011111100101110001101110011",
      "010001111101100101001001011000"
  );

  constant LMATRIX : T_LMATRIX := (
    (
      x"a34051a3a9068b364e3a35e0dd307841",
      x"512eb2d4944dd850ac817c1af5dc39cb",
      x"08dd95491a7f9955b792375440a3b312",
      x"e52f9b98e0a099725d9c8422a05b6dc8",
      x"a937747d1740d63e21cd4706965513a3",
      x"54489933cceadebc5c90d39a754c3ae3",
      x"cd49a4fab4a42339f451d8a6f6e563b5",
      x"61a9abeb8f6b1c988f95d917cb67c28c",
      x"f7626abcbc1fa1374cf4c20d88658b9f",
      x"4c30501459aee9dd4f58d514f8441a13",
      x"fbedd7673621dbdf35e07437437b972e",
      x"81fec42738f2838340c50adcbf8a7f02",
      x"c71a5cf70643258cb12d72721dc29210",
      x"c5a0a3ceb5fce9c165cea64a3e25f62f",
      x"9cc465c0461984888482fe3f0c45aed9",
      x"e8316beaecb34a44be0bbe71d93883cc",
      x"96a562c9cdc2a8304bded55cbada03c3",
      x"a7809854d1640f2859bda1271550e413",
      x"1bb30d5f6658e9f421d660e252a9cf31",
      x"7a61dbe3cd0d88dd664dc3080178dc1c",
      x"57eeec1972f1406ee613468453d0d9a7",
      x"3591f34156944a5bd10e67081cfd1717",
      x"cddfcf49e29057ac2d2a3d26381a4743",
      x"ddb8ab247f4471d69ae1d4e3468cdb94",
      x"d9faa33c5c336c83ca4465b244514ee5",
      x"dd8fef9e19b269e1a28d0e1013ce1390",
      x"2a4fd40ace60db390ffc57e5983444ad",
      x"681853ce04c2a879f02d0383afc64337",
      x"cd51ae395e833f0740f934bcd10642a7",
      x"934efb77d666c3112eba3ea9aa17f1fc",
      x"b73e2f6c9a652eba0f0317db855891e3",
      x"fcb524671f4a1ba2313d46065d6c9636",
      x"fb1cab45b96fa8de966e24bec4e733df",
      x"ad1c1f2f3076c43fd4bc38fd22fd8413",
      x"2e06b70f1e19a9c6ecab056570555c72",
      x"687535530a7bb72b5b16d0a418fc461c",
      x"c208c07776d23eae08766d61a84137cb",
      x"48c545fdd907a602a99bb9c77b1265f0",
      x"e5845cae9b8beb202a56dd9cf87a3cad",
      x"6988cb83cc8773ec2bac30b6f1468adf",
      x"4d537a97f4aa15515e67d9711f2f7fdb",
      x"e983ef05c55a4f6870b8bad0e3ac20a9",
      x"1b44d15f0cdc18ac41e8890934946b97",
      x"332806fcb577f0942b17dece1cae15dc",
      x"2628782c8aa93d86d0e7c35342ee0aac",
      x"708c7c185a17994d3f0877bb419b42b6",
      x"de9d2ec2bc2cfa8221456047b8624351",
      x"74a9b900d20a016751ae2ec266995eb0",
      x"6cce80495102065ff38537c10baac2fb",
      x"fb876cc425e4752a6690b165bfef2076",
      x"724628a023920f9bfaa2ddd9ed2fa557",
      x"8aa2d7b576b2b0b4e0b96afba344e936",
      x"e1e558cb6d74cf0236678a78a212f943",
      x"e1a744eddff12a7ec38075223842614f",
      x"4aa032d8005d49ce98892c73d9d21b98",
      x"048f7ea6fe2a0aaef136da047154e282",
      x"316fd41310e7c7e5c09ade69d7dc2efe",
      x"4bf11f496d63a55d6b3312645476f525",
      x"ca2c51283734fdd501636c86314f108d",
      x"0a888ae95455e2aad5aab95fa2ee0dd9",
      x"e4381ca42fbd296f3a86f8e6cf76ce7d",
      x"fa357b39bbb7d4b1ed99248dbfef1a4e",
      x"e6eb95df50336d2dd7b91179e8c04495",
      x"b3a7e4dfe2239ab6926bc0b41474a45f",
      x"5f53e45d31438675eecf736affc84e49",
      x"9985ccd9af30b166fbcad48597c41932",
      x"3b5ab98696be20d509b5f7f39f37ca59",
      x"e2625964f16ecbb7d0b916b050a1d40b",
      x"ab35dcdaf2da67372442e800fb3f5eaa",
      x"053b73762eb17750fbd1453a131657c7",
      x"b193cd987a16e4385e2a965e8c4591ed",
      x"99d8b2b982fc4718db2fe5934fbc9174",
      x"744eee531a16c078db82ff6aaaea93cc",
      x"9583b4eead8d4880d884d741093a6e5a",
      x"ffc5f20a3844ff97cbfb3adb935bb494",
      x"1b63a0e23aa925c8ee28d0cede07ced1",
      x"9a49169675fbf94bbc2f69e03b781697",
      x"75714a8afe14ef166617e1dbfb2c7465",
      x"32d6cf2272a1cc53aa07b5aad4e71a63",
      x"8fe10386980551830f99994344c3f286",
      x"38de4aec2a19a50912bcb9d2a2e40fe8",
      x"efa95f2fdd5bb4fef00cbfae975900d7",
      x"50a573153ebf76ae576f15e648510efa",
      x"229e02e54f7cef8f2193ca5a6c3fdca8",
      x"3f24cc10ae5dae4545afa9a58088d8ef",
      x"e58cc92494e8d07f22c7af507b54aa6d",
      x"d7bc8879852f74502884a42994bcfea0",
      x"b39558dc8714b24ba07b796e8c85f77c",
      x"b70fd8b2ef9d279602a1d09bc2ab4a03",
      x"bab263b7b85f6dc611d2e44260bbb0d9",
      x"d7d14924c8875db54866058132594df1",
      x"722569ee81185c87baf6acd0727cabeb",
      x"474eac14c6b640ba5f0327e03b4f21e1",
      x"e89afecabbb34d4e577be32dbb10cd2c",
      x"b47c360cf78f35d4615177e075bcaed5",
      x"1bfd4d1cd148fc9c994b1514b7f94458",
      x"2e8092c4fe65b2846fb3b514c6d6628c",
      x"7724bc4ea789d7e5e5baf8872b3aa86b",
      x"1937dfa54e4c9940921f3c5421796692",
      x"34db8057ab9cf82bd4201f4d77dfc788",
      x"28ccbc181802fcd6a04bee0bf11d1092",
      x"8370019947a81d267cf8dcd8dbe40498",
      x"c55678c0770419d7085a4db47c2e8282",
      x"ef273e4ff9afccf13c5d33c7b870e7c1",
      x"e56f68f22b4b3d7755072f3c7634e841",
      x"c3d0839a423beba0c868ae2445a00064",
      x"1502ef5810a21d3f29f50cb19a871365",
      x"cbaddb72abc93466e8195df8e2be5d46",
      x"5d2929dddeeecf48e81306aadec65d52",
      x"5ca1943cd287a8174d38acfc4be8c316",
      x"847901ef1b054de6553eed6a7c794f69",
      x"842b2f82e9bffaae19a5f1fe50b04f17",
      x"5011e94850b95937adb713e74e484eb0",
      x"d43b055f152beb2280ea1bca1590268f",
      x"40060c1b4a981341d743dd1769840799",
      x"975e5a3b184ae8b6c243df5f873209c5",
      x"a007185bc452cca227dbb215f4bc22ba",
      x"125253555245044bda38336b478b2135",
      x"af02fe1bbfd65e178495aef1acdf2cab",
      x"e409e1a6f83592efe0a0e9bde7a424a4",
      x"272da408db6f954af94ade5ee41793e9",
      x"369bc331cebda5cc16a45868497de113",
      x"c3efa04cba7dd140c1e7fafbdc1e8b8e",
      x"c9e751a6ca26f3876524a0423de00fdb",
      x"d988de06b2c89315872227d87584520b",
      x"dbaa0b3e7b49c3d0c8083c23f4c3b19f",
      x"b036e34f9f1dc42e677c3e22b91d96e7",
      x"5719802cf5c3053e782ad32fdd3aef3c"
    ),
    (
      x"cfafb26ba789d1e082361cbd4d0852da",
      x"0034f50ef87832f25cc6fcf1dff0aea0",
      x"8d25f2a98085f192a410099e6f1246f8",
      x"bd9ab431280a02c4ebea15abf335d801",
      x"929928c8bf5dd16662d90e0ec9b22866",
      x"e1ef0959fe4fa117e5f770738d560b01",
      x"3cf80f5bdde869db681f9510318fe8ac",
      x"4be46231a80e5df942cdfe1bc33a9488",
      x"9aef91e9d0bc3618a2602e6d14dd8723",
      x"c446c223751b971804977866ccfdb2d5",
      x"f5c5a08e7190e3cc3c42f8f0839af37e",
      x"80346ccd9ce8f54465a928ccc800feba",
      x"8779071435cc472c66537505256bbf92",
      x"4625721633cde2419ff34f4545b8a3ff",
      x"68e8aae4e0d1ab88e4256b5ca019017e",
      x"837a1a16b16db58b418513567e56f92b",
      x"4cd5b2b905c053a4b2ad4d4f945c9112",
      x"22b5e2772ac112273de1fd80b3095284",
      x"4a784a1d400ba30c3adf83a1bda9bd78",
      x"2696de97d9a609231fe6a827272fc469",
      x"5c7379244426f1dd6e7c59adc5f74696",
      x"c9ee882b04bf09cce039e1d97decf2f0",
      x"f6fc9188f0898857564fdb03d3e6d539",
      x"11f7cf0085e0e616d50b1d8d70a1139a",
      x"af42d4bc717153576994b452f3eb613a",
      x"150e0ddfeca74b5f979d307c563521e7",
      x"239caba64c029353596c7123130f1ae5",
      x"43cdcb00e0b91e936110212eeeafe4b7",
      x"18ada80829b50e92bac3f29fbf8fe3b4",
      x"8cca09177c924bd1006b4b7142e4c061",
      x"5e0c27ad1bc86478661853b763fa3769",
      x"de21c9ae669c7b7167c8a2452b9d960c",
      x"7a8b76fd4dc450de54b298314d329926",
      x"362c940937c94e8a159d09c18dd0822c",
      x"0fb01411a316e3cf0692cfade6e419f1",
      x"b27a7e18b8e60add0cef3a2a289997a0",
      x"33237793e38ca07d86744e1678e6f91e",
      x"e3d5f465ce229791106f1d2d45db06ea",
      x"0413807a2e9865621c3260cf531c203d",
      x"d83df49d065337fc144ffd2a91a9c157",
      x"152c372728d788b4400d6d0fc1b8ab0f",
      x"d4b6735668e268aaa131deee5758b434",
      x"d4bcdb2dd9e9e7ee089885d2515104e0",
      x"52e313c5240d33a95a9825505f67d7ac",
      x"58a16eea0eab9375c1dab5eb826dc6ec",
      x"eee382f9bd248d7baddc8b0a35d38e3b",
      x"693ede1c107756b5fec0202f3a25c052",
      x"c8aae666c932f8f12e31d0c4b088e87d",
      x"be4455567816da21b8739c1d1c2ff033",
      x"33764f63e7fc07c87b1bb68e1f21b63f",
      x"e8c65396738ed60eca2bc8fed8e879cc",
      x"46f28d802b28fbde6c9cb972e5b2353a",
      x"b7bbb47a8d03f66d8942f859554c96ab",
      x"252e863ecdf3195d15436d4afd578353",
      x"13f9049d21a5ee753acf31ff1db86288",
      x"8a6161b75c6c32c1178907333c4097f1",
      x"e4e1633908747464b8a6120f08793a0d",
      x"6eb54cd0fe8b2e9cee9bbd21bf49cce2",
      x"887366b9abe16f9128bc0a77774140e8",
      x"df2e59af2ca9b1dab80175163c0a5e06",
      x"05cf68c6d6d251462ae5d0ea88585e4e",
      x"5b38a874a90d50e2dc06860a98830f6b",
      x"93464e601f0a2c6c3d7d246623649866",
      x"636ff7f1dd4bc9c2620c5e840a571090",
      x"40f7069983a6453f620e5e17216a2ea3",
      x"d6ef40e755f91ef207c356107b1bc0cd",
      x"aaf59efd51bafd29e004fd559029d003",
      x"9af89ae1ad95af450acb8284953de5b6",
      x"d6850b979b0ed4923735678921ed1c00",
      x"c7d643db04ddf1b32d618bf0ab6c2169",
      x"e2d7a48c5b67746115911009aff706cb",
      x"3b99a10bd8c53ac4d237f32cfb2f784c",
      x"5869f4a847a9df808283e73d3af0c6b5",
      x"1a8da57f27a7f5ca823394a85a3bf190",
      x"68879c36db796b85e159d8d420762b29",
      x"b5863b15acf8f9856726c4c3153ffb95",
      x"3514c11bc6bcc9e6134cdd801bbd841f",
      x"9f86c9094f0ff35a60f16ddb4d941469",
      x"87eae5a3ba1d49326c2f6477794ee529",
      x"4c310ffde836e805b092b937296fab00",
      x"b500faee7829fba147ac80d580597c93",
      x"3b6af05ce1673ca0f6ca14e3c41a7c0b",
      x"a552d056368a1919927f196c3e322bce",
      x"4460f59f7cc0cb7e6453c4c2d200d0cb",
      x"031ad3ee19d4fa107b52ef9a21f6b1ac",
      x"1a3b5c943a2bd6595b10b52a24ba1c25",
      x"d68714b0b47a586361d7da0d12a2ca8a",
      x"b24aa365c6c0eeb067dfa6c42ded065e",
      x"e1dcf43d303e20e9734136aaa5957837",
      x"7a63b3a21d27a0300a53a5bd7c52c94f",
      x"ae354fb21f0efb4ed6a36374c2c836e4",
      x"3caff05d8e9e999b5e06c47f2d1dbd33",
      x"19d2e8c3a2d76d01614e72f4ba4fc97b",
      x"761b3988f70aad175d9345f4c6e3ac9f",
      x"136e58a74ab6dbab45c0ded253a1b9fc",
      x"47f63c2ca12cfbaac9ffbf0a5e26f552",
      x"23df74260714764ac28b7cbbaa0e8713",
      x"1b90a07d68ad18354d2ae538996f91be",
      x"f161866dc55223431fd1dea6f8d6db24",
      x"a63d99dedaa540aabc4c2b8743dffeb1",
      x"c9260cc848196473797f6d06284c2e4b",
      x"84500195f5b7218f4d3a677a3bae2ef1",
      x"84dcb0cf982b9148812d73ff43377115",
      x"c89dbe75c698d2b3e8aa73e3830b3264",
      x"a24cad5852e5fb37ae5ad66f90018f8a",
      x"a21dad88aed51b44a2247fd64ed60107",
      x"9312dd81cb64c850aafa43de69a1ec5d",
      x"e2f874fc0b6291436e352006c33e9f0e",
      x"388d9e9a66731e24ceafb2ea6d38d9d3",
      x"197cb4e9e6fa2d2f47ef101d8a087d6a",
      x"7527ff9e15ba40d1bbdd98c88fb13502",
      x"f4035d0f8f65be5ba7420c7a07efd9c6",
      x"ace224dafe58cdb4fa15cf248df7bf6f",
      x"12f9b307217b42f3cbe2220fd2d3229d",
      x"3b54a1fe2a0e0e691f511b7acae3a0ec",
      x"4a09fe4afcb4a2266c0aad2acfdf2c5e",
      x"53c29f96981dd113b1fc99cbc779e398",
      x"2132f5025fb0c17e5ffdf6b618b5c40a",
      x"87961a1c50001fc50719ae2e61191b4d",
      x"90b348cdd194ee1308a68813af58ead3",
      x"ccc840fdd007d771b61ec733930c817d",
      x"35a2996693bf5df6bbd00d789bdc56ee",
      x"46c5381f445b89673cc1abaa4df78498",
      x"0aa108b9e981eaa3c2178841b65ffc76",
      x"ea5f83fc2eb7d2969cccc2d200a0ff4a",
      x"2d621965cdb2fb550417e6875da60ce8",
      x"387aaf09d63ffb8b8027f19e5f15a3cc",
      x"52d47a6adbcd915cb18cef09cdfab372"
    ),
    (
      x"1826cd3d068c419d5069dc36307831a0",
      x"5020fec16839f5e8e2c01b9291702589",
      x"e271d2dd9a73c0e9e2607bbe5c64481c",
      x"1fc6f9775f13ff0bbdf909fdbb31e424",
      x"2615a30ccb7b0ef25e56e2d561f8e778",
      x"cf72d29fa3285e0a964f765dba2280ca",
      x"d4b2e780b88ad36cc80a7a9977fed01b",
      x"06e615ee7e7dab12ceb0ea948a9a2b4a",
      x"9b794ac2688e70fe88dc2524167d58ce",
      x"92078b88e7f3a730ef487f42737be5d9",
      x"94bbc894835571c73d98bf8dbdbb65aa",
      x"63e903b4f284ed9fd7d76a31c4afb436",
      x"714e7f2d347d077b2e84241d01de39a5",
      x"fd57fd3d73ba46f43fd4d34466922a62",
      x"267fa6d6d96932b71979e25aef2b33e7",
      x"f8e7f4918c3f0b49ec881afccb733f14",
      x"33299771a17166125879b5fa2c795943",
      x"c45dfd0c248e2cf0e1d930834fb54f66",
      x"a54168a4d3d3fa3cf0381bdb2be15af0",
      x"b713e0866c60fab63a85549abd0ce508",
      x"fda469d5f765986dec2a39c35ea0435a",
      x"c2340626d40d5e51b978c16792eb522a",
      x"0795fa5b1829745743f1c27fa7236516",
      x"4541a58e95829700f309c78b75ac1cda",
      x"a4a66242d463533431b054401264f2bd",
      x"34552e9cfc091f6bec10dc0ed564f5b4",
      x"9d9b6a2949329d44a1914d7516ff1cc1",
      x"d74a8ef0bd1eae073c011c1d53646d30",
      x"c0824499d2527f25d59f80f2d4c5a143",
      x"0e8f8479455eaf8a12ce9e36942f63e2",
      x"0e51a71a336076ca4a6e61cfca35fb30",
      x"46cd26e0d032b016f15ab41f811f0a26",
      x"3d2ac89f078906a685a7368861fe8806",
      x"98c6473ad53306c21e259d695badb8bf",
      x"16b01eb5d7123da4cd1947b109518f58",
      x"41499310ff3c14a117c183e04d4b06a1",
      x"0060c6d1a42e9ecc35d75a3f9bc9d685",
      x"4f970204b7bb5178f73e5a5765bff950",
      x"e98f56bac7db9e576fde470ace249ffa",
      x"989a6235b7906b289ecadff87d7339de",
      x"ca883fd984132b756d753df643316237",
      x"010314bb4f86474212610d7ee31f557c",
      x"dd4fc547b6d5b78ef6f871a57bc3fb9f",
      x"92771b84c3b3adbafab84e0ca010f81d",
      x"3e55ffb2df889b57107efa94a6c229f7",
      x"5520614e2ab1c6f943a28dcfa2cac2c3",
      x"f8e048c9da81ed5958b92794956b3832",
      x"a969d02f2bea6f9e03fd414bc9519b5d",
      x"2beacd8f6b49a78cf75b58211b1be791",
      x"fbbd449e4ec2e0f9e8979296f4a50852",
      x"6df70b3511d3512b9a791affec45c228",
      x"157a6271eb27a087b370252300aea24c",
      x"64f0a107c4fa3d0c5db62c347adce273",
      x"01d0d9b3f74e89a40cff1bde20a6f3e4",
      x"6af369e8d0b56df118d4f5378acf634b",
      x"c1949aa09e89870b415a8b6489c45317",
      x"fba8bd21f9e64b155015f8707f6f6fcf",
      x"4e2354dd73ea97b7b0f90e9f65e95536",
      x"eeef1e7228a05a6c78f4e48837a1b2b5",
      x"19ec7555ecdbff2ee8ec8c502dfa2798",
      x"493a63b1a51989ece558e032e4cc18d7",
      x"cb2acad84d321ba9d5ce98b1de722eec",
      x"2da101f3037b839893d1a3b0c34f5575",
      x"9b025f80d01584deca2939a6eef24d37",
      x"b8522738a2633d4ac486bcfb14e272a6",
      x"c4d16214c336507811bbfdae84771f59",
      x"5b9a793da12e9592ebd9f578d158bc18",
      x"628a29601d28c33d3196df753b2c449b",
      x"a5ab13f175dfbe3b82acad1575bce4b0",
      x"bfdd8411283b9d9f8dc3638c3a432af9",
      x"945702f15a69504412c4f7b10d6be4e8",
      x"b6bf58f4874ee1cfaff1475c63efd6fc",
      x"c17f392d0f092ebe999556f08973a3b8",
      x"749a87b9fccf4b80bbeed6ee1c674803",
      x"928ef1b827740f37595bce08970ed540",
      x"7f6fff9343b55e253bf9cdc232ea0ce4",
      x"cfcda06655636c515013647372e6a8e8",
      x"d02d5c2faa3c00a5f6d8b7d847ddbf00",
      x"3bbe9cd29ab918a873e754f8483b8136",
      x"65073b6ff7872e0aeb6f4ad7ca5cc541",
      x"41217e9b2405a6dfd4b1ea8411071ddb",
      x"eb6d8f2590e6cd739dd51744360d58dd",
      x"dbcb8b46c9b4ac78e1d903f3966655e6",
      x"076e796033d4a4af62248c2aaaa33cc3",
      x"760cb43a734647ee52f540c770715e76",
      x"a1bb9fb424246e610e9c3c71146b7399",
      x"5d513650408bb729473d23bc1656871b",
      x"66db6f214209e55d46e866f5775da4d3",
      x"7d93c979d3217e868e7dcd096951a37d",
      x"591e3772c43e724e42b9d72ba4fa05c7",
      x"04a336add1a9b98fdf2d18fbea07bbef",
      x"dcf479d2a4f836c819f0759c33e2ed81",
      x"e98f8f1083b22c677143c66263a47349",
      x"f3fc99b39c69302c3988c2f964ad929e",
      x"13766a96b01fe9bf8b29248153abd12d",
      x"0c455e3ae4449fccaf90e8b5af785248",
      x"0382de6f07bfb00822e0e2a47c6de9d1",
      x"b5558d6510d8d89a8baac94b612c0919",
      x"4a13d4f530dab89a80ecf3e3d5b76316",
      x"1e8d327a7355547865748e2eeff3c5b0",
      x"7120a6f70de299823b02bc73651f8608",
      x"5e837e89d3e0ccd6fe48cbeea813d5ca",
      x"d9265efb410c261c5a36991968659197",
      x"296b69eee876174a3e41431c0e791f30",
      x"b85ace62d0a86c6b8eb76b935c94311e",
      x"dc2014352c38f6bc96e627615459c030",
      x"59ef42d8f978de24dc3808dacbefc07b",
      x"d178cc4cbe960f491ec3792f42ab9339",
      x"9b562d04e72c3fe3238e72c53d581096",
      x"cc5c2d01a8ca90f699ea0f29566709c6",
      x"6ae16a7f511c58b6cb4ff8683ae4c574",
      x"305eb0e7aa61251e63a4a00c93ae9f5d",
      x"b19ece20497210a666a4c2b6eef7031b",
      x"34e0c5e076b52f6c265a15de2fa3d621",
      x"0f69ae92b89902f0dee22a2dd5ebdee1",
      x"01512df6ecd5471821a8b38c288941b7",
      x"ee2c082dc91eb978165e82737c8e5340",
      x"75641a96d0626d8fe30d928c9ac2b00d",
      x"659b9055e6fb27bea41a995ba75764c4",
      x"cd59e76648488d897501d8a281dd55f2",
      x"11c5187bb9d2fa9b809e0eb1d90bb027",
      x"db54c702c469612ce5ed019e780f02f6",
      x"e3a69a12d3f8616d115166f3a038a097",
      x"0d7319867b25666af41593b6819fb699",
      x"b6fd486ac71a88d1da62b7c9acdeb24d",
      x"e52ccad214623c6e2d682c78f2f1cd40",
      x"1955b98785254c84355b9ce817c4f093",
      x"8f9a36517219dc9b39452753973f3fc5"
    ),
    (
      x"fb9a4262ed33b5149e4086c576778500",
      x"3bd7c21f9a733b5860204706180795e2",
      x"229805dd4094b071441ceef4bac34c73",
      x"2b1f724b10c1168bf6a08ca9a6226db0",
      x"1bb912c0010759a093c504c199ddce5c",
      x"c2f1810cdc9b2a2b432f44a44439e6f5",
      x"6e54c5852ca5ef14a2f95c19caf597b6",
      x"04b85bfda5c0edcb1e479ce570a20568",
      x"018974358492f3e30526d6b3f1864407",
      x"5dc7f9e037f1e56002b2afd28210821c",
      x"4b14a7dfa23bb91e5342b5ba834a3716",
      x"70ac4778c71be03b7af72af7abb23b57",
      x"ad6e6845ce9e5e4b359de8d6328f1f39",
      x"cfcfdb881c9013e6cb0d4db59171b89f",
      x"ce6be93ec516e53f4245a7fc3783637f",
      x"71b9614553889bd792f8d624bbb09ba5",
      x"5e15e98991566a12608e61bb46a57d47",
      x"c40bfe9ca9b8a819bf7fa3f21df36612",
      x"e1bda98850b35c64fe2615ae46fe5589",
      x"bea8acdde05fad1b1265cc149cc71d81",
      x"95fa3f1b8b24ff6078031de0cc582725",
      x"6643ff9cd6a035f7e7e2f86af0651d9e",
      x"1a6b62c8ad81c9e5f5790a5e734af766",
      x"7059a217f642284c0b7700521063fbc4",
      x"8ee2dae904b50468227dbef07b78606d",
      x"e629fd005aa8c37c9ff55763289275c5",
      x"2e331eec31553d4f3b6cdde2ee7abc9b",
      x"7f35531617ed90d9c0e8b3d228a07375",
      x"c2c93d5ad3f5f6202407c4a8a258f076",
      x"72054be45e615289553919b6e9542ea2",
      x"afeede0b7e4527066650c392d4a46757",
      x"96338709b3a0d325bd25e3afeaaa0cc5",
      x"eebc11614607dfbef5604cce78046624",
      x"c3a8ca9ffcd6876760a10c7fd35a6a38",
      x"267955708693ee225025997aeef73ea2",
      x"52b903b2fc4b7e08b148a6afb7e651ee",
      x"390dbffa7d3031e5510e5636557b97e5",
      x"abcf564dc7603fe205f16d0e900a9f4d",
      x"ba5ae7a2b629d55c97f215ff4f11094f",
      x"a4a90e5353ed5792a821bf1301b03c8f",
      x"9bfa02da911c0d409a946e75fd703cf5",
      x"2786fc16a86be2ee996d2d8b0b716195",
      x"507fa230425d9341871f4bcdca06c49f",
      x"25a5da8abebde3ba762e76bea633932b",
      x"372d8f41fd94e8862ce5427722ba4508",
      x"e336d4e37457d691faee794aec0a4387",
      x"eb723bd0c85e120260a4e927830ac91d",
      x"abb9a6a7620957486d742b870d15d611",
      x"9a392259585e5c61dc5b7fd4ba189488",
      x"b8e2af4b00a295f755b700c36fd840aa",
      x"1ac493c1b8bc14b3dbcb254537ea4bd8",
      x"bc6fd5eb2e676b2d3e675d0e0026a451",
      x"3d4a344be9a53c5c5b354d24800a450d",
      x"52db02df9543a5363df2b5bada72e724",
      x"4a0aed9b0bb8dd5d521f37ba397a607f",
      x"2ef4c1be9ff9571d784b5ab1dfe32b13",
      x"20a160b7656883e402b2d8667bf71fee",
      x"81cd3e85d3b17dda405bc402ab3c5ea9",
      x"718cbc5da20af2e0c0bf11740c7d432f",
      x"9e33215f545d970d5ec0871027ecd52c",
      x"b62914f67c45f865cafba4ca5aa62760",
      x"583c3fdbdeca95605fd2c21345e1e221",
      x"9b4bbf1557d09676a0bba8bd13410b3d",
      x"592eca5287e120f13bcaf5676ac7d4a4",
      x"3d5a16af92192737144eba9af3d3c42e",
      x"0db01480949fd450383c9a9988cb69f3",
      x"e7a1524806d09ed504b75770b02fdcfc",
      x"2ce7af4c7640c42d8ac3f86e8debd0ac",
      x"a415aec40f53b0b0a50f8f6a584a9958",
      x"9db62a5dccd3b6c5c62146ba9dab83d5",
      x"a4a5275e0cde8327322cbc9206395c42",
      x"4601107124a74ac419132ed441de59c9",
      x"ad7468e01e8c5e576a7d8bb9e60755b9",
      x"c70e3d25e88a5dda896e4792e2c6c33a",
      x"24c01f6cce2aec441a72ffe305d8495c",
      x"ae114bac871ace9aef836d843d90b7c0",
      x"a52a9640cccc8162382d615c2b0cdc1c",
      x"39570ee0b3780bed8ab5a90a9bbcfd27",
      x"e79f42469caf7a36974c945c64f5d57b",
      x"c75467f40a68070cb413cc74d47635b3",
      x"22e315be834ee4145134fa8da6e6b448",
      x"f910da3be720afc49dda5c7ffa4bb29c",
      x"a040b13c00e5a8e7a116647b87143508",
      x"5fc61a8fc844898ead5e454a9619c34e",
      x"870c79710cc535cf0fe80f93b61ee459",
      x"7755c75eb3f8fd3bc464aabfd869c438",
      x"a15dd8bd08ba2e1e063b47c5b18b7bcb",
      x"961b311b968c1adca3786795841e73bc",
      x"dd4027b9fb486f39d4ca2b35ad410aac",
      x"3c28104185d43e8746a900cb7b6e61f9",
      x"4c6ccbce4d15864e0302465771f89ada",
      x"3f859720418bbf0a3061440e44efafd8",
      x"4fb647611ca7d904319956685f8a7730",
      x"49c91a1ca58fdde296c11aac4abfd264",
      x"4ad6bd146b43bec3a960b23284f2e0c5",
      x"8fe8364800e9efc5d8a7d3ab5cc996af",
      x"4726dafa7e6b5434a94ef99421a1aa99",
      x"f2933a4f85601a86e0d14d6b164a2a6a",
      x"3d9757cb9d3d02398f625879bf919b13",
      x"9e42c2568f5791175db2986c960be756",
      x"7e4c5b40a60c6127ee6ae99eb69b3ae7",
      x"c4e4fcf4391e4ee4e02419f990a3b087",
      x"ba93f90f62e3f428fff9fc279d2ba7ce",
      x"bd58f3ef11c468b6a762ce131560fb7e",
      x"3cc9841bd0bd5299b9b6f035035a290f",
      x"712bd13117d36b6a0e77f15efbc3320c",
      x"f37bc4a1fce1539d18d680fe502b8bec",
      x"e339919edf6b40c177feebe803da1e70",
      x"032c19186b16c4b84021106ff1c23a64",
      x"3fa740cf6fc9123128992e50b0445a8f",
      x"9c7d4891b36275a86cf021fe1d7fefcd",
      x"20c680d8bac06ed26a1325200f8f29af",
      x"489dcb8f7e7221045b80c59e227736d4",
      x"b8e8219e870e35fa13d0e95342690b6a",
      x"da178bbdb9684e5ca82f6b4988e14d3b",
      x"ebbdc5794da5eb5d3b489f24975d544d",
      x"5da20f9bf92eb6694a923c2934d13f91",
      x"99df2e44411ccc1f577d844af3e7f0f0",
      x"851bc4b62d6640fb145055eeaeecba99",
      x"4127d64130133454f1ca0467764171e5",
      x"0a1380f3e1bda9b387898d2afc7c8cbc",
      x"9b09dd1af9d2bf0c7addac4fe5f8ae55",
      x"3fd1599af63e5a7bb1eb29928828d49b",
      x"459fff15be041f3a93cf2aa0d63c4506",
      x"5c833de847ed181d66e826d47932c4f2",
      x"b86bccd46e6749c7c04347e3dcfc05d0",
      x"f72395b51ec7490308ed7f8f609972f5",
      x"2f251c9563e584f3b0782cac166c9000"
    ),
    (
      x"b6efe08ffe83211da15df5ad7bee9552",
      x"398b8506a8d2edbeecc15d00c5f829e8",
      x"622dc44f79f973baea4d5675ed473e52",
      x"3d773053c1395bc7f3d6b9f94136aadb",
      x"5b310b253aed1665c3ff81c048be0c05",
      x"54530664fc22efe620e3d53792651c02",
      x"f34f9323eed823f5e3e0e73d9ae7902e",
      x"0cd119b9176b2696a0defe93e5dcb045",
      x"27ac59e2e934f0f056f2289f3b20ce50",
      x"2c2633cc2bb205c93ff04332b6e6e369",
      x"c78ca305264a38e6948b3e5097f54938",
      x"3b720fc0b239316d84d76f3ad01d6c5b",
      x"2b4c13ca57ae6bff560a275200fce6d2",
      x"705aab1b5821436caabed9d4587d0578",
      x"eb4370515fe3c50133d05bea8b9a396f",
      x"86512689e267e5ecd7f1e35b69395400",
      x"16a6e2945dd8e5a184962465d0bfc333",
      x"8619afe830c04c6e4bee2279be65eb0a",
      x"bd9f47faf506a543bf6aa46c159220aa",
      x"5be5b3ef44c051088cf3dd283c85b11b",
      x"9f6985a95d808f4a652c3c38f861936d",
      x"239cc6611cdfdac7471d2b60a28d3c46",
      x"5c9ef889e00186b9c6413d3c3f3d4cfd",
      x"a9f9a3b2a517119432bdd6877c8b7585",
      x"8e40e8f21b7d8eaba7baea256a657bd4",
      x"3e32567872fa2564ebb2732e6e6e12a7",
      x"5ba0502eaecab6f778bcdfe85b2add8a",
      x"964a34da07c963f30a0638f3f7c0862e",
      x"c0eac0b51f3c2f5d96f6596005c1edda",
      x"21cf5552431e58d7b69189bfea69a0b0",
      x"d79538328159687e9dbad5882c1fab90",
      x"da40596ea7ed85134433594765d089a5",
      x"2aaccd8e587c0f8f89928f1a42733dba",
      x"d822a426853717517bbce714c38f0a90",
      x"c66cd084b15a40b4b0c2b911f1c1c9d3",
      x"9c0895f80477855907e60018ee2b23a1",
      x"65e7c6879d1bb0d0b9c49bfa32200e29",
      x"24a4d40d06fa930dcce2c23ed563552c",
      x"2defe631bdbd8f02c35161318e1d9294",
      x"ff2c4abb2a525d1045ecaa076f47d484",
      x"45c02b1e0bd6738d283cc4563d0f1d23",
      x"af620926341fac07f4c6618097471944",
      x"9ea1e228c664392ae977419c26cbe9c1",
      x"4b90938c3c04e19868a0b728fb7c1787",
      x"25ac49cf4046ef3fa1d9dc11083a8fc7",
      x"3ced056caab01b95f2b0bc4109ef86b1",
      x"bf0413bd196930856ad73e6e4fd1a43d",
      x"08e42e380fd9b28ea3f483cce1a5aad4",
      x"82f6398ed3360de8a4a802d301624136",
      x"db00f845648552223c7fa8dfe291a59f",
      x"abc6a8b7e0f2520497ba1e958c823e93",
      x"26b8edade2dfabffd9dceaa1e680f143",
      x"5fd09fffc3d76a53c059dd46bdf6c19c",
      x"b4f8fbee3ae2b69c3bf1a3c7f932e700",
      x"f2cede24fcbf6044a7dc069b3cdb26c0",
      x"303b3de55c9cfe2391bbab4c3aae6a98",
      x"4a6262b69e1c2e6f19073d4562586d2d",
      x"bf0904ce081e2af4448008c888a3854b",
      x"b134493a8f3ab69dccec73d2b8cad53c",
      x"26c22504d4ed020c07f77643b7fb9658",
      x"e8d643e4803902e431008456dbad3fd9",
      x"b2e84e0729883a02078a2f5eaff2e539",
      x"64aa30209caee8ee642a8bf62cae5609",
      x"4ce13f73c603b1d94b98efdcd24c5d69",
      x"dc216ed15fc2e07c1b2c045a6fa82698",
      x"68c3dc570e655fdf1aaec50020b53a38",
      x"c1ecc041604bfcc20454f366e33d2c11",
      x"403d7a3b274704006ec1cc5406665801",
      x"b25d9c82177acb54ba7d1068f31a98ac",
      x"fd4122806c59897ef4f78a7a877b8460",
      x"bc533977a44f38fdcb3aa4fc7a2d75a0",
      x"0369f0719d69c577b1317fd689680873",
      x"7ebb9dbca8d2b079c78f82e671687e1a",
      x"94b1c9038be88784e6188db39876977e",
      x"a3983dde7e091527f2673a26b55ec37a",
      x"a9d59855342e17e780640b2b6cb3128c",
      x"45fdcc7e883ceacf69827cd4cad01671",
      x"c8c33a34d12f752498fa588708391434",
      x"9cc0678ba1fad157d8f59a3ded1b9643",
      x"9477802562a0b22a309a1fdef08447d6",
      x"aa6ad1fa54c315dbf5b96ce785aed713",
      x"d01abbc605a16316d9c4ce572a7d267b",
      x"fe8b7aa0d6fcde9b94e2b050cc717bdd",
      x"5d1b532017bf13f2e0b347852f41e54e",
      x"2744ba4836f2007db70665536430ddcb",
      x"feea5a7dcafe09b47394505eba8c20a4",
      x"56c231a6d4f26c39180774044a5325f1",
      x"0a0b5e8cce29eaa0b6bac7b8d9221ac8",
      x"6a672e4f24640b5a8ff2588bcc7543aa",
      x"1e21fc93ce46a9f1b9a7524dd75268ee",
      x"0f727b461f5228b20f560e42631e3ea3",
      x"51a6210996c9db881f829a523da7febb",
      x"2aec1df8fa166e33d65b4e96f4da3992",
      x"ea3cd5b214b7dc184624564199bac270",
      x"7d714b503d408bef3f8ac120886e55b5",
      x"b241307e7eceda998a33995a6de8047b",
      x"d8cc0fc00275119eb02758e77f002764",
      x"e0a42dc5f86acca78d591a47a97c31a4",
      x"b5117632d30391acec1aa41e2ae5cd91",
      x"9963fdbb89e7eda1e96fca871a2e0d9f",
      x"c9d1f3dbd6d1d3decba2ab753d895e6a",
      x"8950f37855b8f8c6180dc2bac9b3fdb5",
      x"bd489105e6521b18dadae3258e655caa",
      x"d46ecdd41e40caa8f45e8241cd795868",
      x"3d2e14e4f231028f467ebcdd8001af10",
      x"b8eed0fa6aae0fadab757984edd2c4b7",
      x"35365fbd930c9acdb4f7e5b58c329983",
      x"3dc48d8a46524731d8f0e65b4b2ab6c1",
      x"f2e5144b8bf04f171e9b0548a5f8dfad",
      x"724d53aec930c0aa238efb75cbafa393",
      x"40b80d5ab21103f096d1b92d0a38fe51",
      x"12f9fac995f2b8b8113d429bb2291238",
      x"5cb892330c359a96c504be22b37e65e5",
      x"ca0fd233134fb01d7f66d8c548b8aebf",
      x"a095cc907e7de30f0353c33da5471d59",
      x"63b37a069a8641e1eef5e5a8cb4ac424",
      x"4695b3c80f8870db8853f5365de6c25a",
      x"32fdac4b2ddbf3888e8e8356bd7e145c",
      x"d1fd84208442ef057c8499ab984c8f9a",
      x"1d76b2678284aef83a70df59bc8102cc",
      x"6795aa2dfcfb4d899f3285ceca27dabb",
      x"e2eef6e2e7f6b308304987c6478634a8",
      x"97a8cf137a4ff64d258159efadd2eaea",
      x"f999d61ec2402a7bebf1f7b96aaa73df",
      x"0328106f22ebb372f89a97669f04abcd",
      x"6f7a49a82b0877872625507367c502f3",
      x"fbc096dd54cd82f310cfe9f0f2407493",
      x"c56d52793958fcfbe25d63f6f102473c"
    ),
    (
      x"381964a883c74c165a842abd1b4208bb",
      x"bdc098137dc90340a074dd069d15dd4b",
      x"734af8db19c2cf11abe376c02674cc21",
      x"9b579965a4fb26681590a82e062b563f",
      x"8aa9b28e1868c49367eff0dfd2652811",
      x"c6542b9d7d9478b1e1cc17bdf95fd83b",
      x"51997ce826a258d49c00b442a42c3059",
      x"e4a96142f0816a35bc0604ceeccc5929",
      x"1bc1b838dbf77f7ef92b4ccbe8440b84",
      x"e4546a7cf91de2cc8d8b89c66b6443cd",
      x"b1decbd761e30cd796e847bc062ddf87",
      x"f2814336a3f9922d7c4b8bb764bf588c",
      x"d19b2c681e40e7e3f38fb2ad04cefbb5",
      x"24e37f0f150e7dc771b0991a8336bf31",
      x"f82db6d9741634623f915f711c53015c",
      x"2a74b1ff10ef9bc158c2d7eca864ca53",
      x"a99f3e25192ba6629358dbe187ace498",
      x"a47c0a38a1522aa69494ccba73425ddf",
      x"4895c8a71b0b9efe63051a83da01b168",
      x"935082624bf876bf61d4df396c16bc24",
      x"20cc41b0e95af63648e324e670596b87",
      x"f52bb9a5278a4fc54870906c66de029e",
      x"dae07aaac783c5b5a6440566f2435e41",
      x"18c185aeb83dfe78c4f1e3def5bbde29",
      x"ea96be77dd0b621ca0c5f1282bba91ab",
      x"1e074b96d7a87602679ff162edf93c43",
      x"97722ffb5e225475356eff49fae5f4a8",
      x"1b2f5c1d0ccf55872c24c6020c35077d",
      x"4c33db78eac5a101f6ef98cfb6a54a7d",
      x"477854510720bf941849dffa2bf029c5",
      x"3b27fab76f7bc23d7ffb8a2ffb4b3308",
      x"a25df7ee539bc4eb3cab8ba71f1cd488",
      x"14590e6c7022d4c066ef0a5963e01ed7",
      x"4e72ace12880947ae127ed7403adf3e5",
      x"43b75800eda8e604cadf699d356e11ec",
      x"4be71e0fe96b6519785def3bf4af63cd",
      x"c1bde44502194e941573913553d93488",
      x"cbbbff3cdf11b06d78817db27c620656",
      x"44eaadc5ba7c1213e7a358391c5f7243",
      x"8303e19bcd6d7e659d010baedd52b10d",
      x"4e4b700f90acb455872eab5f2fac9a1b",
      x"1f2292dec3736600d263cf76d1c2bb22",
      x"6541e02c068d5bcc39c94307e95131ab",
      x"403894183d8db1f00b473bd67f717f86",
      x"92c5795cbeb65b98d45b1847b64b631f",
      x"2f43f757816ee5795b821387ca0fcad1",
      x"fd9f6afb7ff264e569c50b71710db1f5",
      x"b8029d3b3987bef30a1f4bd96dc21b6d",
      x"9f15bc3712152dee9558b7955ab0582d",
      x"27e4c00a1e9b51b9e42de2acc16a2b06",
      x"d2ec0019d68ae5fe037d0eaef3779cd8",
      x"b64786932a5289c7b4b2d134f49ad4bb",
      x"8c82ef203d2c0c799fc92f3ed831735f",
      x"6fb0f2b7c04076a30198448c4cd6a5d1",
      x"0c56aa21f49bd668a87eb527705e3b93",
      x"b86ef7acbf1e6a2ec7718c9902036893",
      x"d4020986397f2d95e17c14ed0113c576",
      x"a40df98465e966d5257800f01af44986",
      x"02dbd63306ea633a743ff4b6b5f946d8",
      x"1f1847ddc0eee1d0bbd01d8639d78ea0",
      x"3d99bece440f7e3b065a0477794d2c8a",
      x"c90ffba16f137c79893ebfec06feffec",
      x"ee8c0b93a982bc0e66d238221627d136",
      x"9a1de538291b56bae48917544fa683b3",
      x"039e07428d0550b961c663b66e563216",
      x"5fbb3f9bf27bfe53ffb95f79452c7777",
      x"7d896c3067a6ed4e5395389256ee3c7f",
      x"dfe5a2b091dd3faeb266c182bbcb999d",
      x"081de2f26bdbfe029b4db6d2fb552fbb",
      x"cf32776fce4be3c0f751aba69b37a3f4",
      x"5aa1d2924e4bb416993146f3315bd98e",
      x"1abf6e03e299849a09d2a38d581a3f9b",
      x"19617a67dddd279418ca8c7528e8de84",
      x"0af1ffac1fefc7f3919ca283a8dd09fb",
      x"8030ed44475d6a8bc745f2e6f2ea8580",
      x"98df8a76a60aa4e9c340fbc48f72b148",
      x"3103d9846502166be3576a730bdf4669",
      x"a47c602d25879deab1c82b996da506e5",
      x"e9d28483b62345922debd93ca0989087",
      x"4e5daf680e414f975c5017dad227a063",
      x"ac473b35df8d55d89ede0806c75a48fb",
      x"ed13410ab5041ce6bc65a249672d288e",
      x"435cf4cb99147f5523ea7b466dbcd3e4",
      x"f1f4d95fc595577caa05ae2687dc2e98",
      x"4ff4b200012bb899f6506df1b39ebcd3",
      x"94a399e1843784b29efdad773ed29afa",
      x"11c561abc1ddb114d74bea56199cc8f1",
      x"f102690eb5db03b93e2b9b75ad81cfd2",
      x"a7fcc48da6484c9845c829e252998581",
      x"80c7c23b2653955509872f6282ba3c42",
      x"dc7347319ec3f86927792c21677d74d3",
      x"df709d65a43dfacf600a20a2142a6749",
      x"d5a913087312f9a2fe5a412282af0fd3",
      x"f632de62c5fd1e42ad6ed7dc06eb97a6",
      x"7db7d92a9a01b8e4536221874acd2962",
      x"430e12ae83d64a73cc7ef48d27a1b235",
      x"e60a5b1c9081e7533233f8a34fa1ba23",
      x"9ab45ef7d9bf355666abf7f7a612226e",
      x"12b082154ffbdcf7eac9f2f2fe857174",
      x"d59be01c441c90b20815fbd25ff1c058",
      x"a785fb8a67443ff55e02c85fecea630e",
      x"c54e719318465f3a4b52c27d7a74ccc5",
      x"4d99a8e2dec319293e6c6f3cf95465b2",
      x"e24bc0b3743907115b7497e85e814e08",
      x"458194f4be4f33f92c788932fc100934",
      x"c9c78ad718b831dc80ba506a00ed1a0a",
      x"5e77a58b0417d4ee994591abd87ff56d",
      x"4b8842dded309b6610c9b2085c6f35e5",
      x"0400fc74e326a5e97037d4a59f67a36f",
      x"d63b7e835db27cb4f1ddda94f94161ea",
      x"74d6d4127c7d7b7a94866f5c9fb7167b",
      x"6ea27f1ba30aebec07adc0d1fcaa8d79",
      x"9c3f4ff559c7ada0427bd49145dff51d",
      x"d37b2bdb605c8c018694b2b6f5d30e6e",
      x"acf89f0d01a0e393d25778fd9ff55d44",
      x"2a7bd68f362ea55136adfbf7e79cbcb1",
      x"0931894bd379264b2d9bd00f8adf2b01",
      x"a5319fdae60d44a0873bdfec2611f04f",
      x"954f7174ee9c1fca4e6633085035e6bd",
      x"07ca3019a84614a45527ea99e1bb812e",
      x"ceb2a00fe3538b4af4d3680e3c7c5ed6",
      x"f83abbad6ac074e0f86a26e71fde5038",
      x"e6f1f1fd7b6b36af011c523345745219",
      x"500f9de49053446d3894011cc642047f",
      x"7ab041bcbc6a8a11a5fcd90e68845d36",
      x"991d18abf58977b133d27f458d3683ca",
      x"80f1d55ab4c27712e68a17b838da92c4",
      x"4eec324f5cc0464ae83706ce8f1ba322"
    ),
    (
      x"b5b81b5a4dbf36f0dc8617c030e0d395",
      x"b7d02f3a7e8e65eaf6ab5dfaff966b49",
      x"b3a88a4100c7b23e95cc0b896840040d",
      x"338ec68133f0de58ec3cf04befaab267",
      x"b42db6831a765c49846811fd53da83cc",
      x"d7e07e7760b05a87dbc8d9bb19f243e5",
      x"4f7c0120fe8c6d9f991892f239077801",
      x"32f903594c7779b4270bda2bca2bddc2",
      x"5aa004157fba57d96ee64e25992c1193",
      x"01a26c20f95251f68cbcfcd1bcd20875",
      x"c6876abef3ca9ac0fec73554fa0f6806",
      x"bf91dc8e99b49a97fc211febc2d45665",
      x"861eb36f1c1f25e2d270e216109075a7",
      x"de177d4d9353e922b888ef8b09b2378d",
      x"9418c58c3b15db452a8e490ed530831a",
      x"675b45ad7564f291b741654bf0833457",
      x"9828866f0ff8c4e40e182a8c1e81e12b",
      x"da9e421a873019936bdf4e66cd1c6afa",
      x"4cd35a6a5c2f162cefb784501061c517",
      x"0c845f1285b4fa75a8a2104b4ccfee53",
      x"27a27e1ba97979824c95e364ac71f761",
      x"a705580088b470209224485dc589eb53",
      x"69f2b499ebc6fc647e40e72fdcd0856d",
      x"59e483d03698c58cdf7e161a8bf3bd23",
      x"c16e8e2119a7431fd43808060624f37f",
      x"75c8e0f0af10b61a24b0dccdc631b9cc",
      x"7d0ef43090874747ff1f155a434c851a",
      x"52b66c030d9f0036f2299ea39bc33484",
      x"9b6ffe3f6c7ff55f4ef157c581941b3e",
      x"92aa1a65aa817eab1b0035b31ca1594b",
      x"3fd93e945d90ba737419f3bbd86fde4a",
      x"035456a429df2486a4275f995e6f3100",
      x"47e87c08797c48b7e2f93a8f6dc064a2",
      x"7b27ee272a88d4a10bb5ead41c8d12af",
      x"da334a8cc56cf5f23d5a58c19450238b",
      x"8e03c0c192a2c304a1eb056959b31e2b",
      x"f865ca068846cc45df6c93a612cf9071",
      x"0b4bde7901cac966f5f03ba83a4992a8",
      x"29b350ba9e75e578b518dc0359ff463f",
      x"79ed003bade8006e7ea717dde8bfebfb",
      x"35db0acc0355d77b9e0c52fb7964b0c8",
      x"e872c0b8929252262ec1f68225491512",
      x"8e071663fdbd6685f6207bd1dad0f054",
      x"8ecff4afbc9fa9e96444936e9aea190d",
      x"53616c0ed8a1d55bbec9e84b75fa1f73",
      x"694bc52dbec10e5f011074916613bf89",
      x"2ed852d23531d6525233599e3cddf287",
      x"155f59c2c44105780b214c54bffcf512",
      x"f7ae509b2b55fe57bf66bb504a8c34e4",
      x"6ed7acecbb396d93549a0349ec0527bb",
      x"566ee6f25303b2c120cce28296651314",
      x"5a525297effd500a3b2a4786fb08edcf",
      x"6465666724526e7d09f6f1b91bed955b",
      x"3f25b36faf34a5150cde2e1a9631cd33",
      x"2be6870378247a18d510af33855dd69b",
      x"9f1c7cfb13e0639667fe5e96dfe30531",
      x"03b3b320b9a3c41ea4d2625064936d14",
      x"32cf3bd291d3f46346b1be52c058f683",
      x"7dc4fd85bf787631b5e0e6efff4074dd",
      x"8537d22f9b9df25c9126ba17c4674814",
      x"c9f826f11d108efb7ca1e3939bee694a",
      x"482f4e1071f1098694b692b4cf3658bd",
      x"c471ba47889f57f483c34354c7e0fd65",
      x"04988a676191943f4f29e6aa3dd744ee",
      x"17db8412b2b0a9027fd96be72fb50caa",
      x"0b2a14bec01bf852cbea3d890b819497",
      x"39da5f8b524f546995b7faed294cb6ab",
      x"e8e54fe7075a8d423b1ab495bbe96bca",
      x"867338b4461925791a8b09c790abaeb3",
      x"d8e6cec6954f1d910c971af5fea23137",
      x"ff3fbc943f6e90c205b71230b3697371",
      x"583cdda06721379f55247ff07b284e6e",
      x"977246b816c2e75bdc2150e401ea1217",
      x"9995838a0571f5af1628b7b500353baa",
      x"190a45849c9a8c9f4470a61ebb6101d0",
      x"23206d8b97fad2f482af060d63ee1b05",
      x"dd1e747475feb8aa342a4e1834ba08d1",
      x"4b704e726368fa523fe00dd2ebbbfabb",
      x"5c041e3593034c795352d4249f4fbdde",
      x"bc6adceba4cde7c30bb692e0fcd35819",
      x"f7f0e668430ff90fd99abbd8a032d182",
      x"c9e99c5ff2b221844cddeade72e58eff",
      x"83aca340a0b08febfef89dd81a6d013d",
      x"45c55f33a604b48f3fc4504bc6f88c5a",
      x"ee9f36873b2e4ca548196ec7ee7e25d5",
      x"27bf0a6904816de27b81bf495700bdce",
      x"0fe02e57b72072452b44a1a42030c187",
      x"b75463d1addfe3d6aad2dbc55ca62cb0",
      x"ca140533e88808b70b8b7723fa89631f",
      x"e1c0bf6ee6ac3a68ca028a2634a954fb",
      x"e509b0b5f57bbf59dd916de6cb44cc10",
      x"5268866596d6ec20bc4f326b9aae3580",
      x"4a2d8db2a0c67376437ba3050649fd0d",
      x"00dbffb3b4023ca05f8f8de8562fd6e7",
      x"e481fcc9cacb546ec87eb328532501e5",
      x"7d6289cdf768f49f6bb99badfc34570f",
      x"f9ea665dac6b516667b0f91426f4e41f",
      x"5f795ffff2c4e768afb4275e53fe7f76",
      x"1b47cbfaedd9f8a2271d9587028164ad",
      x"4e94d35c4596f96899082d7ca97caad1",
      x"118853498acec629627ab8a7b0f2d634",
      x"85ec5a82d363d0c94766a47e4312bd6e",
      x"5de53051a917c7b9ae419ee3e3dd7a50",
      x"c7f56947fe68f23db4d283ac2109c0d4",
      x"8c6a2f93a9844c70fe33a00fb72d7e83",
      x"7e5960602e07f30c3b82e30cbca15a8d",
      x"4c101541ccc8e4f307ca97fc40903e97",
      x"e2da04bc3995a8a50aba89206592e148",
      x"69e6db4491bb02538a06902ec81f1b2e",
      x"77c0f082585f5c5ac3565f94d0162017",
      x"280e2ce73e162cbd52e23e27154cea65",
      x"09ed5e7cf21362f3b3a9e201b2d9785a",
      x"25957e96d117982e2663e42bbe23a41f",
      x"8bf4680f6e5782ed11ed245b70250210",
      x"c6bfb5a9072e6799ad79ba50b572c367",
      x"5dc2c242f41bbcf0679624f3292a45c1",
      x"9957ab77387c13d1cbe88557aec4580d",
      x"2e39b6e40ff91cae2bc6c5c7539d56c6",
      x"01f87fe8ae69f3194d36bebc16c1d6c9",
      x"5c2bbfc7fd11a5c1afe6714a546b6618",
      x"a3e8cb3114d6fd65028399c4e2351495",
      x"5f2e6eef3ee9a6e9c09db666209e89d9",
      x"25062e2635263d567560ccfc82c277d2",
      x"66fa01feb7b7303df6275f0c633c64d4",
      x"e238f9d45ae458a5a4f1d8832cafd8a1",
      x"0d9eef26bc9a04d897af3349fdec4203",
      x"d84434b3538eb32cd2682b5ef29be6c1",
      x"a8b4970bfdea73b241d1e6979e5d6d15"
    ),
    (
      x"3729e1cd3bf0fd33684f0ebf48161462",
      x"7fd964ed659a74de10834404a6e059a3",
      x"91e41d72dc8ec0ff538f8174bb7b8427",
      x"52e05841d4bbadde1f23e2c527569eb4",
      x"9cfe1c93f0676158688a51423bc024ad",
      x"18def7387798823ba30797fe5c1bfb3e",
      x"a62f58c207a33c817c8025a3b6745c76",
      x"f4019deed1a5c5f8eb4bccc9475674e3",
      x"6b592328bca8c9e8cffcdc90b2bb5ba4",
      x"66ed6ad9d8b33e1e77e3a839c1493469",
      x"b69664497f51d3cc27ea507f031c9dc6",
      x"c2e007d3fe80e469080025fca4758a82",
      x"1464b4c4dcecc8635d3f5a87216c02a7",
      x"75137b365731dc8fa79cf2c9d36285ce",
      x"a6bfe7a35669c0b69a8c48b0bba24035",
      x"a37390703baf5185a3509288c15f62fc",
      x"9a80d9417213035fe77e63ad8b549cb2",
      x"569acab19d079cf781e313df8762a77d",
      x"2b54dfafc85bf2f0b3e19f62ff68113b",
      x"d9f0750e13cf075d2f742bee58a454cf",
      x"e6efd42b728534c5211081e38eb459c7",
      x"4f8e10edcb550d9362d87ea3ec262ad0",
      x"d9dc22394d4a15e6e2fcd00718f30ac6",
      x"226aa7c0049890021559f1f399d48a9a",
      x"191cb11a3b92aceb031e7d1dc1ed22da",
      x"5d6ac620b04a9e6263b3531ea27e0c67",
      x"5a64f127b4d9773f40c32e5e4d49a386",
      x"b42d7d36054580d3953517ec6ebe8af5",
      x"3ef1d5bba162d617cee69abc5ce52d0e",
      x"25bf39f37ad7dc77665d8d424caab37e",
      x"cf1007591a7ecde043c557ddafebe37d",
      x"6eaf5031d54225d2c8e174fcfe3fc375",
      x"6fb7c96e7b206853c90683864307640c",
      x"515bdf6a431b4fe77b0579719c3ddd5d",
      x"bbafc5914f6caff44b8c43fd488e767f",
      x"ee178c6791c1ec4bb7bb098748771d90",
      x"70dd4a7564a3d3888c4f73120b160d77",
      x"888dda5d995b01dc723db14d6a680da3",
      x"97afdeabd81c82bc0ce0ab2fb66b1be3",
      x"f03747392615687733be1f5425293763",
      x"49993fe40b28bd852a12b3ca2297a899",
      x"b237c616b3b767d06685d4d825e0bda4",
      x"d980c61e66a06ea5590cce6e3d5ea16a",
      x"6c91f25c40196ad84c3cd91cfd59456c",
      x"c6b0422d20c496234b12434182144d42",
      x"a589844ced91fa6b4588527eb9dde9a6",
      x"4f30d39e61520a124adf9d08e73757a7",
      x"ab09e09bb56f2507ba4a31750e52f0c7",
      x"481d3e77adce966feb46c335bd472117",
      x"1c9a23a2e116ff56814ce5e6120f8a93",
      x"633d078b29244876ab702d69e719184d",
      x"8fc1a8ae64be86a73c284e65014213b5",
      x"13fff1a03ed93429fb43388d962eab4c",
      x"bd5cf9deeb7af3240806d63875f70405",
      x"22505e1587ed252fe87fe4a0fe250841",
      x"f30a835f580136662320f950bfec9cc3",
      x"8b93f1d525b4f99bdcfc2c909465c392",
      x"0e2beada4323e81cbfd690d3341970c8",
      x"168493937df684fbb8a4541082ba9388",
      x"5607c080a4612bc589f71aa05478cddf",
      x"094c1b99e0d1510b3be3e1e74054583b",
      x"cfc04bb398ff17d34b7fba224ff3b08a",
      x"96a02b597e73f54c847b864b377707e9",
      x"adb039c4cf52c68b3d1e591776f3ed63",
      x"ad736ca786f0be13424982d7ae8fc38a",
      x"a6443b5c06f1b4452f1e305f14a23b9e",
      x"8065dda628c852b8ad8c1c567fc2c995",
      x"21005db7654f5b136ba2a357b67d6a2f",
      x"b7d8e3b555d144ca5b9a31e3e4073b40",
      x"b43f678ad6ccb3f694dcbc74fdecc3eb",
      x"7f32795cbcf82389a122c1160bb91a8d",
      x"8d96ec689ba1c43aaa5657edc94cd024",
      x"ebef129fc3139510bd23f3c628ddfe08",
      x"c29cd47120c44d075fa2d37effcce990",
      x"a343b702d63320d43d7963b143bbaf76",
      x"fd18c0541e6465634a9c0183cc1056bc",
      x"3308054326be3baa3b82df53f48e1121",
      x"6ee548691776bbc114e6625e087fa673",
      x"41603a2fb16b0eb61c38d869fd0495d0",
      x"3135436456769098445298c0012359c6",
      x"79d16188e7c96fd72d0ff0c4ff0dbc5d",
      x"0c6b6e7be5ccf318c03442c1577c9ba7",
      x"f5251dcd6262c640124bada7a74ad09a",
      x"a0ab32b0d28adb9b38a86b72dcda759c",
      x"58b09dfd44728f4e24c1433ece3f108b",
      x"3214ca99545789f98d4b69cc95fec652",
      x"c7db663bd0af22ae639e56d2ff5399b0",
      x"916b237d861bcc07ca76ead042a84ecb",
      x"a2093b3ffda55a82ed495a945c84e22b",
      x"80e2b60d119112da5aefc126f9118280",
      x"742ce80cb9f1899ed47ea0ce6abcd57e",
      x"00d770c8a1744d9792c8f9cc3a821ce3",
      x"4940d7828c9a0ca3521f2bb521efdbd3",
      x"cbb9a0136fb87d5786e9d5510125361c",
      x"8e27fffec7a4a773d70b4fc952abdaad",
      x"d8dad665c71ac9ce652118e7f8a14045",
      x"c43aba31de37b8488efcb6a7876c8612",
      x"ff5406829f3868364f38089f48907789",
      x"94a41f0bcd394e3667cbf5e9e3007d88",
      x"344319d63446900eb6039e82364b1314",
      x"764a3303a5e56d5b926434624e2cbe36",
      x"2301aabbb454e87fb3acf8a46a543200",
      x"c0d173663dd2311b5ee77993e3a41a83",
      x"af7ae7f69dbcc392e31e08c105c8ede3",
      x"4aa7cc882c031ade8e89f0eb24c52ac8",
      x"00041095f9214b6144bdba7171b46198",
      x"cb24c52034cad21afd5aec3335851f09",
      x"c2bedde5d9bf614fdbe84b2a9f4e74a4",
      x"1ff378b8a263530b23325ebb5e77ef63",
      x"365b381000ed4ef65573c836f192bc04",
      x"275ca24887ba7a2ac2cc2d77f33350d0",
      x"119957864149981b330d5d5783974daf",
      x"7ca97a39dc5f8eaf0c8f81c697697c94",
      x"4f6307657ce2fe683c4f1ceb6ee99b8a",
      x"099e00c6134c61d173307784fa96ad15",
      x"61d3a76b78b30c4c8cb1c2f88a69196d",
      x"13e15f39f319f4588a8a06e2433517cb",
      x"ac1dd4f07c90ec70eb0bdafc65ce75ac",
      x"62507b25b82794a0261b4216772058e6",
      x"861e18cb7c696fcc10859caa566db8e6",
      x"a91d3e32d0d32dac8ecb0944883c3bef",
      x"0e00d62e10ad1921d67c8021f4de1cbc",
      x"7d852493fc55902e2d7a3ec2fcfbe2f3",
      x"d29c8dd0090be23753d18fd768a402a0",
      x"4eb96835426cc0a78e16e2bcfe5d4850",
      x"f01d38ce4b56c15d87d93f644bdeea5a",
      x"849c84107baf3bd8d09bc8c4b6c6fa30",
      x"7c2482d3a0c29f30d919456ebd463ee4"
    ),
    (
      x"9153ef4de297e6be919fb345de4829c3",
      x"8959c6e0850b18dedfa93178412e4f12",
      x"ca7e7d563d41579f9f24c09acda96f94",
      x"318d58c6dc41380c06fd688e02b7ed5f",
      x"ad6abb2d1795823f47e5eb3169424c32",
      x"7934f362f19132dc80d4d398645fa59f",
      x"4859ac62c1872aa3a0dcb6b481bf9d83",
      x"c79fb6755970a596172eca170b3403f0",
      x"d7c580dc03e7a1d2d9a0e47bc64f7e9d",
      x"8ea1424c5fc412034752600ba750feaa",
      x"8b1084ad7a131f90723483b39db14f49",
      x"a89b8881017945b4b44d4e120554bade",
      x"533cf149c7e8cc9c8594472a82b9812f",
      x"cd6e5c1d57e7bfd7f63ec260aeffb5e8",
      x"aeb43ef5e4f1bfa019675589b4fc52df",
      x"8b9e425653ee08b44b9ec3857419b70a",
      x"66dbbe3b5b4103907f04b487a47db7f1",
      x"c9cc2b9dacf070d0e725c30881201c7d",
      x"726da819d284dfb40567886d369bd52c",
      x"f19baacfc776890abcfdbc3c3128db08",
      x"65ccc83136420d9c8e3d63a49ca3d314",
      x"b31b6391b3011045714b44126a70ca46",
      x"ddbc735e58b67380a5f182f452d2b3cb",
      x"99155ec86f74c746d49677e9918f6a85",
      x"6179b4107cd07ae2f472b964c0f76fc5",
      x"bee55be7f6aee3757a16d4482b1fdf27",
      x"7c0184242f3bd71ce80edf64334536ed",
      x"7e393fb3036942f50d8728de2cc33175",
      x"bb2ddd24611d52930c3941e51686d614",
      x"0da0675bebad622df0ff3275c960642a",
      x"43cb7aea844f81572eafd2c082f7d566",
      x"efbf5ce6f8c14271f8d33cc46eca4bab",
      x"fd883ebbebacf701d8d80d212b97d533",
      x"1a7cd3b8db998c398038b5a84e0bcdce",
      x"badb56eed6cf2fd2631e1b906373d6eb",
      x"745f88f6dd6a8c742cce299396f9b5d2",
      x"266130684cbeb699e94b5d449fd41595",
      x"b67eedbdb4873038afcacaccf3634bb9",
      x"d9ae45f71d762aa50867d868ab4a38fa",
      x"f446bf0e285db209441d13e41b07904b",
      x"fdba415323e7e84ef7d587a7eac0f5db",
      x"be32ac4c0a4d1521635b669d97b099ba",
      x"7def07b5b06eb5a8e56313f21bd308bf",
      x"98a09cc59366841c51cbc3d91f18133b",
      x"6f5a35d6aa719c2e90261bc831d7a970",
      x"2c4e3700d11b054c5c39b31b927cd44f",
      x"3c0963ee15951365e264e062b0cc8565",
      x"cca76a4f23f35befa611b673d9ac158d",
      x"1707cc74794740b039646cc02f8799d9",
      x"a84a776260556ef62e176c7528240383",
      x"bea08bc95599ea04a561cb9ed788a36f",
      x"1762b36e65b873dc7cd3349851613498",
      x"7b8c7eb4e33899e521e1023abbcf7802",
      x"3140defa5e83e625adb432064190bf1c",
      x"1e796051bb4b0993353f273d9e3fe14c",
      x"aa0737b0886186f3aa32c14b6be2c868",
      x"5d96f567ed10e5203ad2ca042044cdfb",
      x"2c49beab35c0a21107996b024eb340f2",
      x"0f16e31846a5e67e38814007a8a54679",
      x"d5a9a87a042bc923d4650c5f709d8605",
      x"46e621207d3965d782e4159807b7d66e",
      x"92d0469937cf74edce72937fe0f7d86c",
      x"f3dbf91d43a0886bb1c19331ceda404c",
      x"88d3f4fe7bbe8906c61c23c8ef96b5ca",
      x"1924b482cfd8b80d123d31d81b902dc5",
      x"d85bf82e28c2635f812ea32c897fd97f",
      x"576eb471ab81f5bf463fa3a6ff85221a",
      x"6b2e79cae6c410b15adc8057a7ba84d1",
      x"e36bd4df5f187ed2655db1127f278f6f",
      x"949ac81de82390e17cd040f55efbd32c",
      x"bcdddaecc38174f6f8e188c7e5d3dedd",
      x"3c4df25d01af457720161bdbe5e86215",
      x"7e55f6805e72c4a3e229c7e5aaf0276e",
      x"669a754a8d422610a57d4abd29d98343",
      x"edd185d07b7a8b07c2ce27000781c56c",
      x"d078a51b9259d1467e64b2526613deff",
      x"94b56b2269881202811960847c90e0ef",
      x"3d95a3977b4e20ab7f9a402d441ce64a",
      x"031fe9a4f3df76492974b0fcf4c72a82",
      x"2ccff23e11731271da7c05234da5de63",
      x"984f0cd121fe064a4cf8ec313b5dc5a6",
      x"0ddd04e7584a69a29a12b593f565bb7f",
      x"ac6c1fc58e86f225af84363a9ec045d2",
      x"83e38cc1170031ae5bdae3184b24af96",
      x"5a0c3b7c2ac69526af8103dd429e01ef",
      x"ce60b081a79a928cef3c98786092bfa5",
      x"4e5687c10b1469e1aa9d9517171d1387",
      x"0750475ca81c3bfccf00ee2bb2dacf01",
      x"977f240f3733d5d78405dab500b2908a",
      x"0fdc4ca75cc670d9061dd317b8366e07",
      x"d96abffc65a9a9203499aaf3e31f5bac",
      x"3bbd102a8c8173c73a6f41357c145880",
      x"becde6976f62afb90e7228ca4a637094",
      x"c16fcc22b19c37ceea9e52723fb92ec3",
      x"7f148b6a911bc59eae61ff4332f8d584",
      x"e6c543be04dd599359840c593b141d6e",
      x"0b86c2ca2d549f4127411ac9addc42e5",
      x"3a4c7b816533509d33be1cc28970df83",
      x"c45fbd634034fef43932688b9d281841",
      x"92e5a7dab01336eeaad8f018b7727de1",
      x"11930dd46527236f298cf6f491968fdd",
      x"9cc91433e0f45eb316f43f475d525303",
      x"2254242cfb231b71969171b708ad4fed",
      x"45cea76b0dc7f26fa602987b24fbebef",
      x"6d731c9000dc702b8c026c45232333a3",
      x"f6ebb914f34ba50aef4e32a1ab1fd936",
      x"f8b296b594bd127143ea8cd9f7ab9659",
      x"3cacf11c868401924a92ee472cd23a20",
      x"d0992eef05ca6164eebbbcf9d17d9fc7",
      x"32e37b004d5f1e09c349ffa7c98d4c64",
      x"1678081b96ce123c7050867f96f746eb",
      x"bd0fd8a342690ee828f2160a4a2964f9",
      x"3048dc9f3b17192e026b2334d6a3ee0d",
      x"3f4b99cc1828aa405a5a092cdcc02fd5",
      x"d8e34ba12cfe8f4aaeb0a217267ff9e9",
      x"fc24013081d6289fd2ddd1518e458cdc",
      x"06d5e5969f36044ff404aaeaeaedc2ef",
      x"b6a536caf243ba183613c27c94fbcb1d",
      x"9bf35bc1fc32c552c2be624e96ea017b",
      x"b0dc980d2234ab3720344c641a152be9",
      x"b8a2af5d59b738aa88b08dc5d8911aa8",
      x"5cc35884814c12f3b2768a7384882b2f",
      x"6a9ff1ba7da58ce2cbbb9ccc9910214f",
      x"b3dc51238369e787607bf1cab76247d0",
      x"1c3d49ff3e0eb02ffb306c10d72e74f7",
      x"b8364a8dd868eebd34fcc4462b0f221d",
      x"4b59dae91a865f38808fe348020cb0a5",
      x"25bc7c8e195431a3474e102e0488dc6a"
    ),
    (
      x"4b84ed0fa4f4b7b491cc3e886c994915",
      x"176d22b361b3e66dad12612ca50e678e",
      x"0a2023790a9620858154aaa0673b0320",
      x"e95004d2955f033d8eb69a08114b56bd",
      x"2409a8d10f4ccd71e2b6c826104e0b49",
      x"0ecefbc5895881f1cfe9a66770a8d1b4",
      x"a3e376ebbdaddfa499751bf598fa3f8c",
      x"372a5cc4e685f8690de81efed5bc6d10",
      x"9fa5cee044286a9aa09e7cbc567caa6d",
      x"26f472860d114f61b5fba333d94580d0",
      x"b02a445aedda5fa520a403aea77cf02a",
      x"39fcbdcd78ccf2b136464afd6582a4e2",
      x"255c01ccf12ebf24800f7c02dd741972",
      x"6307ccdb0072729d0c9e9e485120de79",
      x"c4347d5e7fc30ec0cced7c9b7d70f476",
      x"9cc5336620b1f265063a80b3727e93d9",
      x"c7d9d6619be16dd6a4385058f817e281",
      x"c2e11131c339810724f18f8e4c9fd9c7",
      x"917c0a46f084fa06d4f13c60b7c33c02",
      x"40f60d129b464f4f48e9af01f7348d80",
      x"7330372dd29b758b472d30c4f89c5d9c",
      x"265332be33867ed90f4e0d41c8cd3733",
      x"dc09238e2f1d7c5d3b779c0b3d1912cc",
      x"99575ff23c8228a649cf77ca46de3cbf",
      x"42f8a95a02715cd78503938076ee36cf",
      x"fd8ababb5f3778aa8349378640bd6733",
      x"816cdac18c0fbfaaebb4927e65297b7d",
      x"a0a99be5c8f679ed0a077a12d5a22200",
      x"6ab0ec0b03584dc03a6879d2b3abd532",
      x"6831597274111a570ef74f2352fbf2ae",
      x"767c2fc94084654e151b2efd3459ba5c",
      x"defd9944ec496c120c46736d736d61f3",
      x"d43aa11169fbb7a9df592907c2b68c86",
      x"39cbd8ffc5710c39c97aeae720c83d58",
      x"de17941a3f57022adf40e824aeecfab5",
      x"ffa944efc0b1ab9da4c5d10efb7b98dd",
      x"572efe4782364931989e534a219bb8ed",
      x"1d6b66b3ea611d462815395e14f2b49c",
      x"b058e80f8d6d41ef43ec5aa9bc0848dc",
      x"315eaf1a3e054483edbffcce0a45b074",
      x"9697ee89223e3e4837656e6e0724f04c",
      x"927b032d026925b209d8a638ad0a1aa0",
      x"14d19e5950dac8c9f344001f98bdc65e",
      x"81b87b5f5d248c89ff47bfe68024039c",
      x"1447e4e2e700d2482bf23b56a43aa654",
      x"22b825c9e12adc64cd5685fd8044828d",
      x"ef626531e4799012fddb127b9203fc5e",
      x"69fcf8d3a14db7a963fd8d219168607d",
      x"3659edb5ac3ce020a44b25928899808f",
      x"826f0a2dd41309b00e2d74c6fe63d7f9",
      x"72a931d078ed230526c034d5021b3ed0",
      x"446fd495967a47665b160b456d88c64d",
      x"3685f18940962479a50a400ae51ada59",
      x"a99236e51ed18c3911fa103b6a510116",
      x"bb5099283156cdbc363e3edb4cdf3584",
      x"7140893b0f9d5fdd3abf424778237386",
      x"e6fa6eb761a83ea264c88d1f98838cc6",
      x"7178129abc80f664347f1a06bc91658d",
      x"ee593cddfeda254036f583a0f1a1e1de",
      x"cd06b59eff345d942edfd1785cae9daa",
      x"182d18bfd818bf9056f6ffcbdad72652",
      x"f89906671dcebeaeeb62fc4816d1b644",
      x"fe4df24d84e34a7121e55ac9b7267f2e",
      x"55564bccd4c9c02afc699d06e8286a90",
      x"d5008b45753f51084cc2ba52acf7fb50",
      x"eee97b76a9c3afa203a93608b689e053",
      x"683fc9dbd8fb441f76066e0ac6d06613",
      x"5fb92e3196e3b1617ea0b2423a4c7f49",
      x"93ae08f434f744e234df0fde7a4be3d2",
      x"86d44dd03b978083ac1ef30333daff3c",
      x"66170fe119e8cb8f336fe1e50fac5be3",
      x"300e6e98c72f1d9433a1350a6e30763c",
      x"351313ad6303cae388006e3a39776e96",
      x"d1fb4ddf730e3a4f665d82d475fca426",
      x"a4c3d45897bf5d40b9fb512bde2cb0d6",
      x"23f025734aaad09068a99c9b50c76c7c",
      x"b891fa62f67de892eb0515dd3073b3de",
      x"555b7b3a45900b397bfa12fe8989072b",
      x"bde8e41fda5d6148da3e7a0f0ea824d4",
      x"ba15be833cc4c5c62c1b4166af9e32f5",
      x"1928314a0c74e5106aecc80f506275a5",
      x"98ab0388d8187f114285f9e24299471b",
      x"9c6fe678c981471551c3a77ff5798c78",
      x"9b0d8c215685795914536f75d51991ab",
      x"833e3bfaf3d5b19ff64d5a2fbd82258d",
      x"74f5d5e241ee905185c946279d7be33c",
      x"1c1073ccc78293b3cad69f4dd4675f43",
      x"9a13f534900998355b1f045628d07e77",
      x"7605c589de3dbeb5e0bae159a6f1b6a0",
      x"262ccb76e713bdd3d93fe05e62dde193",
      x"daf05f78823127005c69cfc36d39742e",
      x"19268643f3b55c93a4c493e68282e7ad",
      x"a50d892f1f947c3a338255b892f8251c",
      x"1551657cef51495d605f28e60f97b3dd",
      x"db5378eb26acd916c9addd5238f6d81b",
      x"907d4b1f466ada92a893c4275fed104c",
      x"5a29a1835e8ba0ace92a3709acc70edb",
      x"f485b09012646c0b3d9193bf8556e10c",
      x"2dd10105ac62548d57367462bcd34bc5",
      x"d337aec0a2e178a6be77cad9f64a6035",
      x"698b24ffa44c121ee0cc08f1faf8722d",
      x"6a4a93bcf0da0d5103c40d1ccf9b3e5e",
      x"0213896bcd091cbae753b35e137fa2b1",
      x"280a58088be8ffaff90da6d84b3ea198",
      x"9ef214bc38560a9589eb8a386f7530bb",
      x"b91f4deab2acff64585f05865498b12c",
      x"a6358977fb0dcf99d8b9d2bb0861987f",
      x"4b587c3ef9056442eb17fbdf0b9acdd7",
      x"59cda7bebbdfa7d1bce12bd9865b5840",
      x"ffc0006492242d5d29bb9bd6aae33f92",
      x"f5f957f8ad7c09342c23103a6ee9530e",
      x"9c01812085e252d42c7c7a5401eb6c87",
      x"da9d867f7d19c5a84dcdc9684f416bdc",
      x"bedaf2deb846413ce3af9bd2ba5d961c",
      x"41b1329b79e77ff17306cbd6d20b8af4",
      x"92032d2219dd962166dce60910181f60",
      x"4fafe0dbea66337eeb267eac3a85372c",
      x"c0a7c95f9c80839e1836ab85654a0e2f",
      x"67ac9c88419485b578fdf65b5cac1c62",
      x"ebc226df5c7d6c0f9aebbb5cafab341c",
      x"11c82e55b3e576ff9ac57e0cb4887379",
      x"a7e1c876bf7c3f5053e1b8b7e3849989",
      x"f1e5715b649358e1d7f4888481a41588",
      x"f74dd818fecc638bbf224b27b0d23119",
      x"a240a9189da9457ab4c43a1f95758f4c",
      x"811cfefa10cfb3dba2eea61099500865",
      x"9ff4d381a812f66f3d3bc9cf43e51d61",
      x"76e899b32c368f11ebdfd2727a5f3fdd"
    ),
    (
      x"4d40b94d7410784fad69b9967232cc05",
      x"6716bc1936785366dea43ab3c0d188a0",
      x"e87fe3367b71b1da0f7a786efcfc5a6a",
      x"0157b6d6e1e07f6f6d480ed57059c729",
      x"553bdb732405d4b721c855d87732f181",
      x"b3ce5d195b074997e55151bf572dc927",
      x"5eadd16c3f4149493a6ac15c92d7ed0f",
      x"31d9c400bf6f66cd8bc39cddab857859",
      x"4a41d9b27b96a848b82211504c2c4885",
      x"dedf2e7d7bd6c3d419347a4e7dd82980",
      x"2970121d4b9b6ac56c94b2a356653260",
      x"c031df95234e254f3b2f2683b81efc0f",
      x"928ffadf9dd2aafd96944a9f53d21181",
      x"ae58590d8196792f03ba2137b05f174e",
      x"61041131337e362dce27948c01db9d7c",
      x"210b697723ad081bafdc287eacbbb4f5",
      x"a9e637a808888ac899c92cbcd75328b3",
      x"f23ed576a3e0cf1588da6c6ebb8ba59d",
      x"ea79f7db9963133bdafa2fcef541f777",
      x"107868a26e9975c3fa60a2fa4abc41ac",
      x"7d273bda7be25421ead9ae1cc6c86748",
      x"0d085a62e110fe117a2bf8f0359283e3",
      x"2436aa125d087e0a4d29500ce7531e7b",
      x"6c8056cba4f31b6fa8916722c6c67802",
      x"f22e772414868b24befdc8600381710f",
      x"72d04d64d64dbe23ec0633ae4e275773",
      x"90b8acc2d722421f3f69ca5bfea43e26",
      x"38e8b07d9444be524cf420de03f7f5ea",
      x"0ab20fbdb0adf3b82e34f8c1579c1850",
      x"eb02a6ad00044fd70267ba61131dee3e",
      x"599bfa702654110e196217faf230a37b",
      x"66792215518cd10fe3adfb90ad726613",
      x"6e492b371a838589b1b73a018a19439d",
      x"dc699bc57a0464d6299064f941a07102",
      x"2d8e7c5d6d53d6779ea710739431ab01",
      x"079b0741d6097ab1f31f90a3bb62073b",
      x"b5e05ef645e5161f5aa7ce1a8d7d0536",
      x"e82eef94c60c30da8d6a0e987810944f",
      x"1faa9d374d610c6c3b0f8b42c21ac98e",
      x"4d660beffeaaa894f41c55dde56141f4",
      x"069884a09e5eaed023ef14d6d05297cd",
      x"22ba56742347c0703c354c80d11e531c",
      x"a82f12128305496e600c15681e94693d",
      x"6154e3834dfb40e30b591cfc8f76a8e9",
      x"abcc227f595fa7f3c3197b052ca20e6d",
      x"10aa79bc817f18fde88b8bab8e717e41",
      x"2162a356fb4a62fe1446ace1c595bb61",
      x"8e81d2159086bcf4e9501235c6c8aceb",
      x"08a32456e8e1fd417dc1cb6fec7fe0e9",
      x"36417e027095d063d9a5b136aa6bb66e",
      x"291fb930b5c34e44abe88240bed0cef6",
      x"9db4a837d02b06ca9fa5b80d5f716336",
      x"ca79dcddff4d7ed81652632dc959b3a2",
      x"a2b6b6afa66131759859d56ca1e91a7b",
      x"e474b10b2f91be6189647cb8dfca434c",
      x"d66e390dee822ada0cac281b8e0a375f",
      x"a17594acc92b0d0947998227b838f308",
      x"58593273e3c6ae6c822502e125851532",
      x"90d9b8b3ee63d988e17d82403c5de1b2",
      x"2aab4abeb8af194915a0fe7957de6fa9",
      x"1c1db2e64072e7c5f3551258f74bf8d4",
      x"059ba116b1f88fa5441a8428e543ecc4",
      x"5e2edb079270c6aef17861ab208d6857",
      x"7659ba4c4d747af77b9720de7b2fabfe",
      x"9c21a75ac3f65b9d93405b31a43f5175",
      x"0eccca2eca42dec1cd4175107301b0e3",
      x"d74a64eddc3ba1d64cd0854e0022a142",
      x"8f4843a1f0ff10f7d5ce5c0d18d5c544",
      x"c26933cf9f63e5fe1b4c59c1c6c3a0a8",
      x"f83c49ddb593d022a1d5a0ad898e5d6e",
      x"04a5c5e7500c6811d8b4675255d3149a",
      x"f31421cc7ea7221af2842e3c486cb979",
      x"5573e415560e78b4ba75f77af30daa89",
      x"e38af697cd88d8b345529870daf69f28",
      x"a213aa79c0b7f466e9c7d9e4c1b6c811",
      x"aab91dbbe7ff21e29f99539f0bef8f0b",
      x"08879fd0335a72a8c8f66d4d6cd14edf",
      x"06a5e2c9dda64da17393a4dfd53fced2",
      x"59600b1c5f45c0c90d6851d300a1d613",
      x"a76419735a572aa0e7dc3e1b8c524290",
      x"65ae6061e94dbc270b562d09b0ac1b8f",
      x"bd75ca326c839ee2a9f511083abe2b4c",
      x"b7c5882872ab919412ef4fe69cee83aa",
      x"a0ccad79c43c227d294c84e266bb15d8",
      x"314fceb231c8df102f3344fdb8073d4c",
      x"1d54a8efda50f1ff75931bef1ab222c0",
      x"105b3b8996dc33f5d31f8185ac13b133",
      x"c84cbcb14995f93f798474c3eedc3f83",
      x"ef48f257a83ce252838302d9500ce9a4",
      x"53100a0860f5cbc55d5af25d7b4bc440",
      x"e1fde5072bb0598bdc8e4cd6239c211a",
      x"a93fafcd5c86129fd70f33c3e1925974",
      x"59cb52d3824e2daf044b2135650edf89",
      x"04aa5ca34f94c14e94f004d5cb336783",
      x"1a014f9b14bc542d4c55da71055a16b2",
      x"2ef28aec23c20a4e0bf4d1129b4c623c",
      x"44ddc62b2f70b2f0353bd043fa92bc71",
      x"0830b9bed4f802b26619c6c7842bd354",
      x"7b9994134b9e567f3e1c96d00b4c645e",
      x"a509de8de6aa7e000d3f9b1ee2e4e232",
      x"9da7a749f1339de6b32cd918808fe517",
      x"0e13d0cac923b4aec937e8f3a948df64",
      x"b1dcef196603927fd8041315dbd47831",
      x"6ce582c6ea783e71c4b40b65048c826b",
      x"a08ca3001d1ae222cca2ab878a506991",
      x"ed5332e34b959bd1c1e98da8576faa3c",
      x"0537a6d5c14c2071a4b0397c9c368d9f",
      x"791c7d1d72e0762dc96a35db25ccad14",
      x"f79593f3efb8fbeb573a1888e01be507",
      x"ca8790685f115e78c1feccf894e06aff",
      x"f104814e20959b9475d3f776423d7d6f",
      x"cc455a0bca09589be7e0c60f73551255",
      x"5dfac938f8bfa9d6713f11ca07b995b2",
      x"3209fb071e345740c5e3c05ab8f1b809",
      x"7c04080ac95b7189eeb3e43af3f31e99",
      x"fb92d2adc9b11068d34bea9e33d08a2d",
      x"ea86f624bee2ef2eb31b8c97dd9269db",
      x"7522b457a6bbb19fa2fe69ca79d3c84e",
      x"477eb6e0626ba6c3ebe5e1bb2b01d893",
      x"a7ddd024f8fe52013f88f9bf6022fb62",
      x"d61b25b61ec1e6718d34e6d40076bae3",
      x"0b0e54a2e04cfd2cbeb3c29ed1ab0028",
      x"986ca568e664843798ff5b5954f80c39",
      x"64211eaf9bf5f9c19af00d1c3bbd0760",
      x"9534818dd795982047c4e7622ec7828c",
      x"63b34eb5ad0fcf39d75d56efb4f00c0d",
      x"ec4b357ba6107f26e224e8640642eaa9",
      x"edc136ac5d91713ff38c40735ea87a71"
    ),
    (
      x"a01b5789eb84bb3b54f4f594d00e7b88",
      x"aed5093e61a7e4cd1c00c124abca3983",
      x"1d53a0ccfb12304677b111c96e6e50f9",
      x"91b72af920aafe3319ab72425d2bc09b",
      x"fb6565596a9e3a8deeb02cd82e08f549",
      x"fb29a142ed0ab0e6211c823881efb479",
      x"bebcda5c993a597c2c0937c21de04077",
      x"cb00a791cc6d456d058fd9c9235e2b0f",
      x"1dc4ffa95bca1e7881f0698c65180c88",
      x"effcea1530f35ef973983f3fe589462c",
      x"500c03b1d108a8cf4ae08884778ae5b6",
      x"c5fa942871ff4a28641a2c09d45969cc",
      x"64fda203ddf540f6149912828b609574",
      x"a5b566e069557c533c89e6472d858a66",
      x"6c1ea4eeaacd91c065763783aae8c3c9",
      x"3358a109943e34056ace72988d40f19f",
      x"04d08d52b51c56603f0c51cb67a61c6e",
      x"26852df996d00a6da712383ffbb9dfcf",
      x"4324ea04d21086212297e76674756dd5",
      x"c6ed4074075b3e45b6b85e1e5dbc1453",
      x"d07a3d7c4946f78a2bf4927971ce16ae",
      x"170eb003ac505615a1452c50ca0f4e4c",
      x"823f68f7c99a974717f2b589880fd347",
      x"05e606234ccc43ed2ac326c8870ee715",
      x"dcd8c756d2fa66e26e1da80a5fc9485d",
      x"1a1262d0d03035df3d55a80e3ebac656",
      x"76ebfd00c3bbebf6332a0977211e5ea6",
      x"85c8b8ea648784af2558e863d288a37a",
      x"b95301a34f4e6efa8e7ed0b85f365428",
      x"bdc7cafe101bc2018712e3deb72d6106",
      x"ebfd2c5929b0dc1b02f4e9358fa40ae2",
      x"d432cfe697fe725624c988858821a621",
      x"f31180d4c65f0541a9c488f6304ae069",
      x"ff34c4d4545f999426073c95e311f978",
      x"d7623ce4513ce572e94d421d311199df",
      x"b11ea45436fd4f4e0cb7c1ee270b8817",
      x"813ca9e1a0a8320791c48584efdeec38",
      x"2257e4d412b87db7e76a12af9df3e173",
      x"43852c572057d1c38219e5f5b562b902",
      x"a0f3cb58c3cf5d51472f4bc9e04645c7",
      x"303f10ce2e4598877c522023546d647c",
      x"7ee796eb500c9ce765997aa9ceeb7372",
      x"6b25eea77ae7ec7e89e4eaf6c8a77fce",
      x"96b7501692ea5f4f4a1905c77dcb93b1",
      x"64b9dde41a7355719cb7ab8fcd1027dd",
      x"4faf711b9c3c219ef1f548ca426d5236",
      x"08266e7b8e8bcb59ffa4341d5218bf52",
      x"ddf6bbf412f9f1e1271eda81cfd1796e",
      x"eeb28a3372c5cd3d074c136adc2228b6",
      x"db81ab66d7fe134a21f7a85ef40eaa3d",
      x"729082796ddebc1d93d8136946fee9bf",
      x"98392e28c0bc844c9618b6a9c4e665a8",
      x"404839c4593b3fa64e6e05602f55f9f8",
      x"362d29acdb1d1a702dc3a19272284f7c",
      x"ce7e8ff2844efca432dcbbd0a697659f",
      x"21ecbd58eb0a5cb44198f07cad6e3cfd",
      x"6ca03dd7c45555227258ff9929691b7b",
      x"e597f37f506aa27713d22e2d5bbd3ac8",
      x"b69b792eac205fbdbad54e23b07d26a0",
      x"2b16a425c3eab45c04cc8a0bb2285b17",
      x"341de7613209f6bd7294c2dddaa4a51a",
      x"b6adf5094e0915cba6d14ed04a6f9215",
      x"b53251fceb206d2ec8728b78e5359369",
      x"236652d3ddaebb202b51d1dfda5884bf",
      x"eb917262ad33570e2060f523d3266794",
      x"85c8bd6178320e9e67004368b8da68c1",
      x"d66da246021104fe3b97ff66cf68ee4c",
      x"422a2032d3b7b67d1c11dc155629d3a8",
      x"2312913d70d586fb7b15134c20caf7b5",
      x"8964c442e6820f545d2d0cf8f0b9cdfc",
      x"9120f946e54508b344c1bdb9d5ecacdb",
      x"4552e9755f003edd368fb2cddc09277d",
      x"3fe1feb766cce5022f40b257c57ad786",
      x"f940762b5e5ca021b7c2caec2c432593",
      x"04f9d2b44101cf8099ba76e555f8675a",
      x"2a4f79c17fe681197fb034998de633b4",
      x"22c387e52b1a93319361cd983aeebee0",
      x"e975a4e73d100a283d4d2ae3776d3c36",
      x"48ad1563605f89faaecadbe6b41863a3",
      x"ea30da5cd3104b4d1f5ea1fcb6e47de0",
      x"b87aa7923f92fb61077823d4a73fbf16",
      x"01d2442980ed571972d142f20e0d3cef",
      x"fcadee5fcb9025703cee96bf142b2c52",
      x"a5ead2808197e920b50cf1ed1cff7551",
      x"fc4a0ba3c804bacadaafc53a96671016",
      x"69fe1ba1a887df5f8d80d8d5679d284e",
      x"eefefe4d639e77a8ad62b70761a59700",
      x"5b2261d91a3f5eeb5b44f22b88db774b",
      x"92b4394aaa066d5221c4a506be0fb460",
      x"65c8b571bf328b2c9a676cba3aea4037",
      x"508e56590e9aae7a71e2c9fbb73f51fb",
      x"ab6e0e42371a43b8887c4744159af082",
      x"f9789cc84492ccf6b90e51a02f1e864a",
      x"ddb174b96f2adf464a3489f9728f0dca",
      x"9bc2bf7727689935a61a57fa7eaa1f8f",
      x"59dce99880f5c7bb559cc5f62e963439",
      x"aceb63100562f444afd9baae1f18f20c",
      x"5a046ec9b19ca639b94ee7e3e7cd0015",
      x"5e8bd59bf669e685bfedb12fbd6282d8",
      x"aeafe5ee219edda347ec8599c21725ad",
      x"2ddf566fc3ca4e4c706b90404e11b9a0",
      x"8723437835fe4461334f060011e65a6b",
      x"2a141670e8682f7320574707a3e766be",
      x"525d3783e1678924852270beb8a0cf9d",
      x"b952db9e4e9bc626df67e561f6f5bd3f",
      x"07b7bc45ceaaf56bf151b9e8187d43d1",
      x"e82531bf63efb6e9eb401c1e3dd654d2",
      x"10135abd923dc6487876cf17958b09c4",
      x"83a4dac7dfcde6805a5d054122e8b2cc",
      x"edc25c4bf3290cbca289a15f45b04db6",
      x"ed76d9d41b65c5f033178ce79518b4ff",
      x"dafb50cf8295f459d12268f9495407ac",
      x"fb2f0d580a043b47edf46439be91f4bf",
      x"217fcfe673bcbc24d238d0604a4cb16f",
      x"6cfa377e1d16442f6fbaa3bb39cfcdf3",
      x"e0722270d6bd47ea558f1ff0bdde7b5f",
      x"0b13cbf48a765b21881580370ebf6eeb",
      x"69a8ac4ec729b0d4d552335bfea4f1bc",
      x"be78655691f0f6e96b53229dc2f1bfca",
      x"5c86b22fb6a6aaf2928fd5bdcac42a63",
      x"e1c8f7a326cff38b9d2660b02460021c",
      x"25312b43e2e694a2bfb19f9793bb21d7",
      x"41ae15e114237bb999faea60c6590fc3",
      x"f83dc4ebdcce2127f5b879ecf72e8354",
      x"61d8364789da97efa78ff4b3439c5403",
      x"719bd08bd17045a363e071b54fd813b1",
      x"6da878c154429e3a06a33e36d2e0b6e1",
      x"507832468a85088fa290eace43cf8d01"
    ),
    (
      x"322791805ffd955341859158a99c860c",
      x"d891813e253845548254e9e4892a7bde",
      x"03903ea6a5f002fc4066d3bfa2fedd40",
      x"2080bf7ee496a91b228423051f6afe71",
      x"9dd3b100eb58a85811775e778f016314",
      x"1cdabaace563a598db1cd17fded74186",
      x"baf69058bab9e7077b9925e1a154e1c1",
      x"fd1b9f40909140a414ac44c9dee9146a",
      x"707cb18fa358dd56b519a7af56dd4b4a",
      x"a6376f7b55f45df6a3809feb552a0633",
      x"1fee8f960ea2c13b2547188d7b16c901",
      x"c7d60f6f59cb382d304a2e2731efb486",
      x"cd32df461a656206a9efd71e785e3d17",
      x"93d6a87f0d712d1727b0c97f3bbfc248",
      x"3fa7f6ae2824238e75e428b14527dbf6",
      x"f82878680ea44256c6802207f44f5545",
      x"4b81fa3c46c1325d39fbbe4b0acd9418",
      x"f4c6824058e23587210ba97893e6d34e",
      x"ca455f2f0dc1e4096926569e23f5d202",
      x"b220262ca5b295e4e4353f79c0186030",
      x"6c46570a8359cd88d54f9999736c27f7",
      x"1f583474aeb90c43146fb29a11dd68b7",
      x"41b505eda98e7f2b69777e90c1c25877",
      x"b7035deb10ccff3cb8f060be3e7220fd",
      x"e66c9e0f581db681a1062772e8c8ca9d",
      x"a4c613a443cd72e11804d6a938faf921",
      x"6b38a2597583020df66559202941b59d",
      x"34e8039ea83da8fe481d97e66cfe5ee5",
      x"7332c22b0792ccbf0a6ec6099b3f8735",
      x"81d4e97924ee083bce5f79ec07fb31b3",
      x"ab06801ae12794906442125d49f0294a",
      x"260d4e73f42ec2032a0ac6800fa5593d",
      x"6d8240857c1291e99d31c1966a73b4d6",
      x"27a492e5ec3b1e3b0fb6b7d66d87faab",
      x"ddfd6fc60692a760fa2bef2304bbbd9c",
      x"adac3984d33316cdd040dbef66160568",
      x"c1dde6bfa9c1f1b1265a699848f7fb75",
      x"63a1d9cc6198b23ea583114ceb7d360b",
      x"e4aef3a1eaf154bb713ba79f34b5e467",
      x"0e48358443f6f92bf88e28701ee1085d",
      x"f89636519c48752046b72f4b7e682461",
      x"bf69c1f93d3d7b80deae8af228e84248",
      x"2b4908c3cd6a381d351d0ff06b674c8d",
      x"e73e93f0738127498a32f9fdf6eadaf4",
      x"e4849e261c96ca1895fc086981acdb75",
      x"06a27d908b486adda223018f6cc2bcc9",
      x"e6d3e820ba235d70476706a2a80cebce",
      x"74b63107aeb2ee54b5f41fe17f73db92",
      x"298fcdfbb9272fded37a9d8d4c1acb27",
      x"d3debdd1bcbcd1906e5c607597445e26",
      x"4c2a217842925c90bf19e8b8dc327398",
      x"113887126099c14da350822fe406e307",
      x"54fb83fd867e5ac7415526d723e0322b",
      x"5f4781fdbdd90c86897219a740d3855a",
      x"c8e674a8e45f0e9042eff58702fc12c8",
      x"3973d4b7fc470afac63496ba9ba223e3",
      x"26b2348972593edf0785f531aad57dba",
      x"0121257db31c35eaf4da26637c4d4e5f",
      x"419a960d71d5a5afc282211f2870728e",
      x"189c0beacf054dac68f19f97ba2c4c92",
      x"36f5693fac223f1d0efb667d87429add",
      x"0e002b8491ea7e1ed65c580e31d6fab7",
      x"39df199700146723c1aeb99d8b0d6ff1",
      x"83ae8a40ed49befd954bb1b9524b99b6",
      x"2e24c272e01b2352c9eaca4fc6ee22be",
      x"136b971acfeb94552a6bcbbb8512453b",
      x"59a0c5e0f84ef269e94640e8c9602460",
      x"9f73e7f72cad94d92c185fade2e35e0d",
      x"9134c306cab1b647e06087d5f0fea577",
      x"49d0cfb0bd9d0e3f100c2060660d6557",
      x"dfec3fdc0d4becd8c98913c0581841cf",
      x"dfb6b0ed8995117050d11ba101afc388",
      x"3545d261112872449d7bcaa7b573a7d3",
      x"3f58123c3012d743c5b98e033779adbf",
      x"7beca5a15a688eff1ca5ad274f42695d",
      x"c87678284866cd04da5f5dfefc8c8ffe",
      x"7ee7f58bfc0fa0c9787e9ea41e336513",
      x"44f24df1dceaa36445019e769105b73d",
      x"c22f67d0e84ac02f8b616f95a3869fb2",
      x"9d544d373e7d3394837c2b92d0352b4d",
      x"0cf906d851f28ab909e51994a299a6ff",
      x"11558855cbaf1e9d7937c6b2d13c238b",
      x"1600bed949057c85e3dc7676efdc9b8d",
      x"1b8214cad071216cf792aa1dd4622744",
      x"7105cb1d197e449fd0041587e5988964",
      x"e70fe9b8968bd2b84b516febd93dac41",
      x"9356bc8ae5092b756b6226841a32f9a2",
      x"334d1a51ff2b9e1c9b0f54453f5e9404",
      x"c043ca43696b3f703716dc8dcdfa4ec2",
      x"ebbdac0d3066ab5d0fe0bf6e5887fc92",
      x"1a98584c73d92e775ddfa64d63a84b36",
      x"204b34748e4e0960c295ebacaccd87a7",
      x"2913f40dcfbffd1532878a8371007c22",
      x"dac0eb13992105d430a054b94102ba0d",
      x"76c7329ec7783e9374fbab94b117bd6b",
      x"0ac268ade329af10c3b6a63e568a4ed8",
      x"ec3c64876e5af6a23e089eca23442191",
      x"762a6c8d731150ac85d4427cf4220413",
      x"43c602b5ee2c892043b77175f5d9f1ae",
      x"5053187a807c53d595b5b31912be8f3f",
      x"11ac5a3e818a39a2f498f44b8f0513ce",
      x"4c7cf971fd0735e74f5b0c0665aa5a67",
      x"4c2415a5d21a70c4497e52a20a3e9a56",
      x"c053875cb45cc70794735dd5501c1655",
      x"b0987cbf205f31c97cca681d659b4b3b",
      x"092ebab3b678f7a1e4b2a233785550ae",
      x"6ef60ffc776afba513e0f5ce0ca64f19",
      x"0ccdd6948b30c982ab79724bd1c098c9",
      x"072de5827e5f7c4ec3daf6750d9dba69",
      x"99f5114a47e7e3b769dc255c49e6acd3",
      x"f667cb8085b828a61c53d9e56f2eac14",
      x"43b71b4118ffebf6a5737466836090d8",
      x"243f6302a1cb1b429496ef0c2722af82",
      x"272c086fa44e03a3b53e206b7ec45d52",
      x"5efe619c3d82102cb0ce4faabb7e1861",
      x"f5021b071fe174e6e09e0bb2117816f8",
      x"649ebae7522fa9bb8fbde4fcb84242ce",
      x"18627bcc145901bcef2a8810f19d337f",
      x"133bca43bda4d8dde63c6ae86816c225",
      x"d70ed0c5df6f0e987ea4c52dd738ae0f",
      x"cab85906792b30b13146f61e99eeefca",
      x"ecf101cf88993c8aaa6255bfd85f9be9",
      x"c52cf9ff09a7d72c71cfc82b98796ea5",
      x"4399792ce006ff0250ae5df2db79e68f",
      x"2401a10d524bd736d386b2ed2ae36bd8",
      x"c56811b78476f3943fa6a863dcf7e828",
      x"610081f0c4c48c9190fc4ac727ac545e",
      x"b1f2cdf8a7239e379c7f8ac17bbfc766"
    ),
    (
      x"ce1d5fb9549bc925a196cef4290ecb4a",
      x"027bb8ca10b6ef614dc7ba961df3929a",
      x"524b2e13ca3ffe78e5e99a6acf20ceef",
      x"7d77719a32f9cb42bbfeee627c9a02bd",
      x"f6ddba6cdb5fed1e86490ca0f6384f4b",
      x"186627fa6a9b7f649169b9172865b411",
      x"45d5876dea9040f3cc4fd5bb6ebd794f",
      x"43a6661fc789f0ca37ec4f79cac3a5ee",
      x"47aa0fab57edc9c2c3ced5cd6a14ddbf",
      x"63dc871e4612df99634da40d7c6e018c",
      x"66db4a49ba7565e668290c7076d65e69",
      x"ab76d2de5bfa1947bede1a71840a2c99",
      x"3e8c2b5730b205ca9087bcb0ce2d7bff",
      x"3ff5d25db763c71c25d1614623ffa676",
      x"9042b7e174fb7fa3942caa3d7fc3f9a9",
      x"44f17e5fb9771dfe7d52e11ac0bcea97",
      x"d50c4c8bc75fc7a41813994a1a1b5175",
      x"b951ef7631c6d42fedf79523266adedb",
      x"a088ed77d9ef3139ef1237afdacd0fb6",
      x"a2c049131e9da31a4190209c575eac54",
      x"0b4da7f041262f08f199127e93fea50a",
      x"6c000e3073b99b8534ff4d5ec2afee51",
      x"7b4de1910a2be20ebebc7962e27e15fd",
      x"5b6eac4b5b68014ce00c68e8a468d8b4",
      x"353df3fae9d9e221e5fa5b1626010a38",
      x"0f55246fb037fe8b128eceb0fda5c5cb",
      x"8199cff3a716574b2ead05ec06db94b4",
      x"f3ded17ca958d8f8b5fdf1b0e9b4a2bf",
      x"67047dcaf094d546d0e711927ecb280c",
      x"3a509732e06827900023a664d5fd0f65",
      x"e895fbf388b4a8218af0e6e0be344f7c",
      x"eb3edb433ba8a9cbef34f05da8bdf3e2",
      x"bc1e01b28d08a89b914e5202b3fcfc76",
      x"0babf07a688e3e5e05064df3da739765",
      x"c26d4155083d18add1028f34dbcee3dc",
      x"974bbbb3ba2ab0691d0b36f6c12ef864",
      x"c094952e2fb43755d06c0b8e0a436c1b",
      x"049142675ae5f88f9335406381966433",
      x"d6374a4d1872e256efd83a9dc7971575",
      x"ca4e6daa453b73640b7bbf7791a069f2",
      x"c54fcb6040316f51058881fc0e5a7546",
      x"5c6b9bced13fea34175577bd3a7c6cfb",
      x"907c29e014477b51ef5c7183ce055401",
      x"438e703605a894fd4528de452ed85b7a",
      x"62eb45ac879b8bfb1d49f72c3636ffa0",
      x"0060b159c7f37d8be9eaec0c14f38b7a",
      x"3444baaa4535da300dcadeca268aa006",
      x"56db1925ec677d842fefcecb0eeaf5ad",
      x"54aee205da62e5153e93532123711a4a",
      x"d2f1fdf7c162fe58e40d0e3d084403ef",
      x"890f09a7ae8ecf559d2f259ff131af9e",
      x"6694407b22eddb085d8ae3e559805292",
      x"0c0be2a61641a7b502f27738a722956c",
      x"718010734d0d08956911a5cf4753e115",
      x"ee796c6d8586f3d01688b770c5fd4b6f",
      x"aea77a3590644a307899fae6f2b65267",
      x"574aa5bf2a0bc8b11f69c56e0e042ee0",
      x"b573c566d6ca503f6f57a093d230e9b3",
      x"68d9e77655189778b6be4232f3253ccd",
      x"6138861572241ebf65d219a0e39b3267",
      x"242edf54b8ee954c9cdc7f778e12d75e",
      x"87f7e38fd0bd05595d6fbc65d448ab7a",
      x"fd5421c7e00ef34fa1ffaf1c391be50b",
      x"cbf786259f89f4807442c54cd5bfab80",
      x"679ac08c8184a7b5eacb176a55bc3da0",
      x"f6a00c4592199f4adebdf4ba55509374",
      x"faf9b337aa03cd62747d9c0c599304d9",
      x"0c044d132bc23a9addbce8288527d76e",
      x"dcd8a7d3ecef03a911d25ae6d4f0f2da",
      x"4505835ea27415aa8540563b707a5638",
      x"7cd96ece13a4cd6baeccef64472cd1dc",
      x"e0f9d2152db28a6dc8e927b5680fbb1e",
      x"d38c6413fd31af409d0c118300416d27",
      x"a7b189c1779e410eb537ee52526539c4",
      x"dc4d836d2f741f240b34e23ab4b5c16d",
      x"bae30f0589462e6b5b9187b6c1127494",
      x"672a96732c1d0d01af7befac439d1e80",
      x"7ade83f990b2b58c9fcb115322bb7764",
      x"23ae1a46cda763ffb5f67e38ec9dc91f",
      x"88fb47df17d08d7ba7b20d5146416149",
      x"83c87f7362fa28a03e3ee27232400eb9",
      x"01281f1017414a5d24fb0c1353df113d",
      x"aa59eeebea58c345f11d35d4da878d5b",
      x"f9c9e38dbbfe3c53df3cde1fb7a4ce5f",
      x"16e2ceeb8c304f133157d0569ad36fe2",
      x"29e683e4ee95eca3b6bafd682d7e6d91",
      x"4b3d8ac8ecc97342c002dd19a4a6754f",
      x"54a49e4e1cee741f935341aa9928c7dc",
      x"4ded800f50d047268243e8855367ea03",
      x"e1f5a1991a80871852cf765f771d0ca5",
      x"5a9089cd1cc0c1dd35a3dfd88fcc0bd6",
      x"3ccb16b78f8e8247a5448bcae00e4d10",
      x"f3a81bd4d781c396e3625a7858582437",
      x"b7131ac795daaa7c4a02a6a6c8f5c7e4",
      x"0830e10f945f664d367c68ef91ad1bf6",
      x"254e1acdecdd3ebea70d8aab41267ee7",
      x"f30ac42d1e42a6ef182462abf70ba147",
      x"34176c81c7c61f0ab4a9d16ca8b618b7",
      x"a192a8db1914e269bc99b0d0a8a17e9e",
      x"70aaa7d527e17fafa9a8674848d84459",
      x"5bab77cdb0130d895ab9721cb3c1b9c4",
      x"c77fba609ed4638024d9b0a250f4abf7",
      x"3114965ffe7390ceed737c738b51afd6",
      x"a462b94ab14b21cdee1280396beeef40",
      x"f86d18b64d0d00920179ba13510f2b24",
      x"9078c09f21f76d31b24c54a7043ee5fe",
      x"f5aa44b3c897b7494a0e60734d4a44f1",
      x"6635ae2c0e845dd6c67bc45c3aa70155",
      x"9875dc6e90e157b429936247a68ebb5d",
      x"25bbbf81aac0958f51fe1460f8188708",
      x"4b2e1542324f90a0992d6536f15ac149",
      x"2ad453b97c55013af85b8924b366fc26",
      x"bef89486b360b23f0cb6fc6d85129e00",
      x"09e4b3df4f37a2b2e27bc3a3c8071331",
      x"7a26d6fb278fb656b3ee60273d80399b",
      x"ae394e3e8638a343aea1b0c66ad4afb9",
      x"9c6f42af16a62650058d006d0f31c80e",
      x"5402ea8b702c2ad15c74ff286f5ad3eb",
      x"5c05a9721231253d0a67f0f4f96d2024",
      x"63cae681f6eeac7d4a02763142f8e5b2",
      x"1017228cdb56053c02253c77c551f4f6",
      x"b7bcb331907cf35fefd79cdc56657649",
      x"497de275b6c3c22550b9acd94cd52306",
      x"5919c0b960752757c837725db4983e3b",
      x"d173411ec1ac7b29c8a7372c52b9e2a6",
      x"ad1e1b55a08fc48331563d54a9ce36a4",
      x"05af863eb90bd287dacceaa9a5ca47ad",
      x"e5a016f3d8971a696fb68e5c786e0777"
    ),
    (
      x"f1a45c634725323a8c37880254a15449",
      x"a5c132c39ef5385c2ee4ba34931314f7",
      x"f8764d2822b3f748802d476d07ddd990",
      x"675478e8b73ca5f8f6148bf1817294e8",
      x"87d75e2b2873f0ef692325fb497386ee",
      x"c38b7b3cc67a97e66b2c48f1f97baf9f",
      x"e357b3c45fd0b860ed00580f85ebba50",
      x"19570461e0d8c1a6b2aebc9517788572",
      x"9ff8307a76863e05df76439772a19222",
      x"5f5ab861d254a8af789c7f76efaffcb3",
      x"b57dd951b754a9007fb73ff49925ec65",
      x"8b626481b5ab80bd84d7ca5fed1b9437",
      x"24a2f2e8f975813715b01892033352b6",
      x"80ad66ece2c747690236404f45fea7f6",
      x"2659c19a0bfde4cf5bfc9ba47608c473",
      x"c0e245ab7622ba616ecb39c1d6702301",
      x"9c68af6c5f6f4e1769fd5d1499fca941",
      x"9a9acd4aa7a334750c27e0a1801499ab",
      x"38bbc8c6a960fdb708d28e9ee8dfccae",
      x"d7027edb24c0a609361ad7beb188d683",
      x"240132ae5ae28155f1cd683714c176ae",
      x"80d6a7b405df42d09d30ab049cbf545b",
      x"c67fe7f54f229c9737bedff323324147",
      x"9b579ef9207a77ad5fb220c4669de18a",
      x"861afec9a773aa7e4c5152ace3d20e16",
      x"73f3e4b612bd2d76b08813751b79a113",
      x"8ae5d26b941521aff2bd510ec9ae0ff7",
      x"c78fec21a00bff8f05198552d400df77",
      x"42c004727c76c0b72b38fc8b2f64feec",
      x"06fa7584f7b7110a5c9036956d7b0a2e",
      x"686817cedf28cef357dd1a7594fdffc5",
      x"72106053d8b956dd15ee72e1f387f13c",
      x"0279b84a95b4dc9554cfd9cc6856bb09",
      x"c11a8072e99d808ad2eeb1f412894b42",
      x"c3e0df14a01622a0997085a1f9229562",
      x"61316aed531e72d6e154f46ab3877369",
      x"831554ef8e36e0bfe85e579217ea19bf",
      x"dcb33f16c65c2ac5f49b946c2f4dbf1c",
      x"48fc9cdc644375f80229979260134734",
      x"59701ea7be057bf27cc5e8aa1028a733",
      x"b18392a26ddee38bfae29f587655124a",
      x"22a3c4ff520aac7da921d48e61fc6380",
      x"2d4f2d36126028fb7cdbb36fc6f38b64",
      x"cdcf7cac57d62d8ab8084c900b7f34fb",
      x"2fd256971b4bf05a73aa7c866f1419f8",
      x"448c13ea28cb8b099ebcfa3df2665165",
      x"4f48734f2de39929c17da923715422f7",
      x"81e959cb47cd90d5959371c589b73aab",
      x"75ed1dbec6c564bc1aa2ef0933d820d5",
      x"0e527fc4f5fb1c50fff0d4cb7ae10864",
      x"1fc6b330643bc829ed68e3f35ad24fc0",
      x"7d6a954a49c5ac21491f12d317051c43",
      x"bc0a7f2a1864fc1cc03d19457c6d44b8",
      x"86756478e034d266ce3f190b00f95216",
      x"d29a29e800ada80371603421ec677735",
      x"1eda757c854e18e4d714cf8bd26c167a",
      x"ed4ece67284774f2ac6775bb66f050eb",
      x"888264266b0681297aaf741252472a0f",
      x"0e565d682910c2ad48c94d7df262b0d5",
      x"9ec104fa0c8daf9b7465e763a44ea427",
      x"7d42aa278e6a72e37a0d971027c96ad6",
      x"6cc2a675fa197c3bc51e0e77253146d5",
      x"e1d674c04fb00258c982e5c4561bca17",
      x"044347836c2bafb80e2377b77fe455af",
      x"42ff24960bc73924a011ddfaa285b190",
      x"8fc39f28a153e515b677ea1b3e403222",
      x"b9161d1767199d9b3c4c5306a0f0b214",
      x"12c9a54cbab7b0acf2a8dea518673360",
      x"cfad267035326ec8a5c7f466ee63b14e",
      x"41fc3bced33ea4c997a62d74cf0ed2d3",
      x"75557283b1d99bd7a9ece6a2b201ccf9",
      x"4d957afd8f57001bf20694429162015d",
      x"6303e54dfeacc3f1c1aee0aab0ec3424",
      x"508571dc67568f7afba474d4df2c7a5f",
      x"3b994aa7e18743a35bc68aa2855c7221",
      x"2f08ebe535686fa3faf9f0c38770df0e",
      x"c8d844f1a1c152f473f59ff7457ead0c",
      x"5533ae2834d732ca485e2a85f94b4ba2",
      x"b0a6ee9293008e1854f8c87080079e7b",
      x"545c633ebe8205c8c5c5e0a6021af370",
      x"d44a92340046c7c39c4612bd53277585",
      x"e0528f24dc99eb30eb014d9064d0aad3",
      x"ba59f87d22093828b59374cddc7ebea2",
      x"e4f20917e92be6ac6eba926cee4ef591",
      x"bae606767cca980061237f84741dba8a",
      x"a8eafd7d00e0ec592b9730baa162387c",
      x"eac7d5afe20a9a22ee26dca1a456a01d",
      x"6205bb0ed90bcf2e20763cfec26e3af4",
      x"798f0218ffc36b93232a07d27d4a7a2b",
      x"3504fa056a043f1d770aeec184576d58",
      x"c6097f2d6c42ac0eb78f9e717bf0b98d",
      x"5ddbf9330a4b674926399ca44816ead0",
      x"a41b60132d8207073425f87969b56656",
      x"bf2551d32a2aeeb22a2fe4c2d1020a3e",
      x"5d162e9d1704dda689eda5cdcd34bf03",
      x"08deca0afeafd801ebc4f76b00ccba80",
      x"d9e4eed56e18cbae429649d1fc1945c0",
      x"8ff89e68323fbdaf01ac61ee186c9bc0",
      x"5e2e1c70c9318280cc6303458aacf674",
      x"3b11716210564153f5cf8ad115ad74d7",
      x"e4aa2dd7edbd1a6dedf506c97dd22da8",
      x"3eee1848ca1b63c0779b5e3f86997781",
      x"a8f5e63e33fd6fa68b9055e60804d777",
      x"bac34221c9f00c4bc326888ce251310a",
      x"04c55f4fd5a63b8b44c6ff489e5528cc",
      x"c046cba27118199f94964be29237b9b1",
      x"25b426731d4ef1952fc346704abb7f06",
      x"1fa995b6d173dc1c104582ed53e697e1",
      x"c2e42e71d907860a0fa8d423ca009c8d",
      x"00fdd33787b89ab1b4a629d135589f93",
      x"2f32a8cecc645dbc0e7bae0c43acb053",
      x"b1ba18366eefc0cf2d6bfdf890c0d0ba",
      x"b8b9d66119e69b1a063d7c348df41014",
      x"a0ac4e5b89e6567afc912a8f6f158d09",
      x"6a174bcc0fe8b0f8a76ad16a851d9cc0",
      x"7a2f0493ece4249b9a12099aa568854d",
      x"65171b3be6241803c9537f85010563cb",
      x"b83ac3c7848c38da08910b77dd071688",
      x"cd602d1af36cee42f5b8603bc61de56b",
      x"b1537bf7e7b2a5fdc1cbda3c04f048bf",
      x"c6919b90ec7b271c8d41de4f839aefd8",
      x"6c24a4ae866e06e8b0e55db130cdb5fb",
      x"1ac770711f92b1bd5598e93931132375",
      x"76c25e93d88f548c4d9dcf0e5e3003d1",
      x"7ae1e1e29f590fef3ae51b4d405240ef",
      x"c302fbca96875868c70ec70b7e380182",
      x"7e26dc1adbb3fdcd7ff4ff7672b9dfdf",
      x"7feeaf5c336d235ca64aae176efaa388"
    ),
    (
      x"eb48f717e8977f131601eb77b6ffe1a2",
      x"8d991d62a993032a56a55fec9bb14590",
      x"093bacc4d72d3089b5a26f0b60fa16de",
      x"fad8489f901cbe519bb8de311924dd73",
      x"2cc3b75251aeed89e35113eeedc8a91f",
      x"afbd713bbce348c4245a37bfb9b3ae43",
      x"7089b4f1944ea564ed7f02db0910d204",
      x"729ff9643dd9683d1ddb2daf28e4dfc8",
      x"a7dfa3cb7e937d4a9370cfe0e24a107a",
      x"4ff5ea69e0697e2d12d795cee0628e12",
      x"83df562ce6171f5758e6969f948a2762",
      x"8653ffa6dcd592b45491b66efba3b460",
      x"c4187850cf872cf96e3b2bb97bc6f2ad",
      x"813903294e02bbc0572447b1fe5dc266",
      x"e0b6ddec7feebc7554ae330bf77677fe",
      x"ced531bb31e8a5145e22e9bdefed68a5",
      x"c1f4783be28600a14958931d7eefa46d",
      x"53445e7cc7c68dd424d489d473505391",
      x"3ea802a6dd6fc58eb453192572cf094c",
      x"e9d6e0c680c10a12bf08e8d6fdc43cdd",
      x"5393a67aa1eb8e83357690fe4533f6c4",
      x"d75ea8a2fda952b1e27f78113aababa4",
      x"0647c6dca90242ef4b151699fdce91d7",
      x"5e90b7e0fd3be5439b0e3d46fef1b13d",
      x"9e841f144e9c8b31db9a4486c82e1771",
      x"59f724418fc1aab7332ec8ae2a3def3c",
      x"bf659bf22168c762a08835d2779914bf",
      x"c09a8e8ad3d7b06141b4b1525bd5c1ea",
      x"2686c5a1b98c84e1e56615de0d675dce",
      x"ae9c6795c601ea5d585d147fa91111ad",
      x"34577685b20494f71c5959defe2294c5",
      x"f7db374ba2573e5599c8b63d5bc526e5",
      x"c000a5fb1e0bc6db715abc5a21c5f026",
      x"86b3555c2a335301121ce0659d457a82",
      x"7bf18d0758640c37ee864a1a9eb2ac90",
      x"64e357d675ca4327b8ccf51fae632030",
      x"557ed6c54719ffb5f22fcd1fdf2f5769",
      x"9c1264421843ca79051c945f0374ec9b",
      x"0d5bb2e6a603398d121ff88b221f7bcc",
      x"d9696c2d30ba46fdb4b4fbbdc261dd18",
      x"410961b5d220a683cb4152e59d4deb1d",
      x"e58016074650f37f33729ba18612c99d",
      x"70942c05c1cfc0f53fc80b3a5b101256",
      x"b55fc234c867b89e600956939c0c6c29",
      x"80469b2408cea7ab1e1c4686fa21c793",
      x"7e66826380d4b8b2723df9cb0d03450a",
      x"38dfdd772f76c4124b38c88bcee8bbe1",
      x"89408a431161958fc0326974ce877c87",
      x"316a50bdecdd149f12b425229fb1c293",
      x"bb5133d265599f35f28e5b20861799a2",
      x"c984e94aadeba794d1599bfbe60c3ffd",
      x"cafc77de547ce1f9d9b0aeff852f6d17",
      x"282bc7e1f05072cdf2698154e3bd36e1",
      x"95584dcb62527bea7f72f8cfadc5316b",
      x"8b19934a4093ac1e16b11cf34bd9627b",
      x"349545fbb9860e2b26f284db170dcd59",
      x"a275abd731cff4582a550170b821bb08",
      x"851188b0efe443fa14ec1ff8bf66fa9c",
      x"de58a3fdaad9a0c75e6e23909d0d8824",
      x"39dd702f33e70c7dc1f9da46a78c5503",
      x"367fe2248d7aa9d6a21ba18048e96837",
      x"a77f980782417834b8500eee28d62ed8",
      x"377877c87ef0686bf334fbc1d1a3f746",
      x"1b4bd1f76461336d01b3ef2a0b28fe59",
      x"213bf4ffb9db5e18a427b4f021591753",
      x"4606cdfa44e839b8daa1535c51600c5d",
      x"3c56fb53878483efcf2e36fcb4ca9f74",
      x"650f300e7a5b6e4c4bf6fc2a662f1671",
      x"ee00b50edbb10a806c10554dae43e313",
      x"b63ff0853542598acb2c1abd3c57a9db",
      x"92905cd3badde2567d01626977808b0c",
      x"1a5e0304b8f483be84cacf79d90c00b8",
      x"721df7e81bcf752153a164285b8d6942",
      x"d8a8a3cb6bc516d9d8604fec2a5ebe49",
      x"57a68df2d1e23af4e43dade97cca655c",
      x"05f93bb57a7e28ff9a2d5098a8d6d7bc",
      x"47a8933b664a6ec098c811b7f7ebea5f",
      x"9e0df805181d20a87669d3366454b4be",
      x"44842e7c220cd64cc111acec7b5b986a",
      x"547651457cd52fa78c3ef9d2f6824909",
      x"8b404941be2bf23cb8cf33952cc3047b",
      x"b5011e73fc536565df12dfcd5140182a",
      x"8ab7f3d15b6182adff8aa7a3a5f85029",
      x"aae2093488b8b34231e5745e975570b6",
      x"ba8315cbe911a24fa7d39f78494523fe",
      x"e24aab0175ae413a9ed23f7a5f4dfb5d",
      x"e0b94a0e6c3f6a346def7bcb227fb925",
      x"7917116a97287e635c3f0b2c8c726426",
      x"dd00f2f90d2cd3967f13a7fa943f0ff4",
      x"8b567cafb1e75fddd2f115774c12b93f",
      x"8bfc8ace51b7e7e391d1453742d09fd8",
      x"d5ef08fd3bd08d44225d5bea66b9b42f",
      x"3c1aed7939697bd6629a6b4d5589e39b",
      x"5f07d8e46eb7d20daf1c8c330d26df7f",
      x"37215f4d8dd829fdb3a4040340c5ae41",
      x"c044e63d4208e2ae5386b288f8e5c030",
      x"b2f1415e8ceda8f06387312c1fd23969",
      x"449f41ff9ed20562e8e075cf8aacceca",
      x"33a0501b4c4b4064dae8b90de8a4bc75",
      x"c846799d0980ee0439f4b57a6118458d",
      x"23b68b9b433fce7abbfd0317c229910a",
      x"1a4a26550bce68da68637410f10055e8",
      x"560483bcfff081f7377c0776c397b771",
      x"5dbf12ad916ae16cbb4f6534383085cb",
      x"f10d0141e2d7cd556cefddc380ed4949",
      x"0d1538edb58f97d983f12fa5f84c33f5",
      x"2bc93ce2289517cedce99d8ee4ae4ed6",
      x"f27834b77fcfedab6616ffccd0d90346",
      x"863f3520ad19e6c3dcb2d91866389ffb",
      x"384b9ed16a1551500647b3c37690b4bf",
      x"3f49b8207d99653fa3240a7f925aff8c",
      x"fa3fbff721fa1cb9c09f368ae7d621f3",
      x"8198d91e36f3e3de9cdbf594f45c1d2d",
      x"634f84eaa34ab3a2cbe0cd8cd59d3e67",
      x"a5ad7994cb78e2a8c2b266e1bdf6c982",
      x"bc17483a6f88a580ad108009ad8a569a",
      x"48210036b889c63d0b668df50aae9142",
      x"cfaf3b6f3d9afa27ccf60212a4f648c6",
      x"319382be22d73486225f1b03cb53c516",
      x"a63d45534f8a83332b0bf3d46bd5da3c",
      x"759a2e5f55a51fcf6bb05cc122137cd3",
      x"3038953845b60e0ebaf336226634d7f3",
      x"31df182f76141e42666b52f8609e03de",
      x"363702a06eb68e541570125051d21e1e",
      x"8a752de2336bbfb7fb2c11cda365d600",
      x"a8b7e8f9d37add7586a3a7143334f4c5",
      x"00a3f92a74317bfd5c2c4c81d8ce3663",
      x"caec1395bd3cf0a04e0128089d5707df"
    ),
    (
      x"dc2fb38a74314d1cf683f555e3a6be74",
      x"e51d55c9c96738f254fbe8d1936ef452",
      x"faeed1574f5f59a43aa6a9784c84e26f",
      x"b780c0ac434b4a6cdbc3c40f295e6569",
      x"c9ea08b30993a27525342a2bfc7b049e",
      x"9e42db19a0a37748eec6272643a5469f",
      x"966220b009b66a8e787b63af60c75601",
      x"7cf5ff9004d55a17d58eedfef476e2c2",
      x"1196d24165c9ad0105e492cdbbd18b84",
      x"53ba8648aa60e9c27f80200b3594bbb4",
      x"17d91c7974a787ae369a5874c2a88481",
      x"4cd4e599e92e8fade8828c89afcb5d54",
      x"d743a7becf8faf5cefe44d22203b6946",
      x"7d0c53e178f39435a33683d5f06c9b8c",
      x"f6f11485dc9b9838f3f1e5d8ec0ce2f5",
      x"6d10002186422f786559a70d0ca435d4",
      x"18b08fba05dca0b48654815160934f90",
      x"ad0edabdfc91600117b8c4a291abb5c6",
      x"c6a449fdc4eaded7e337f075455e3edf",
      x"b2c4512e0845fadca9a136534e35dd22",
      x"6ba8ce845c1e47f302dfbb011e34fa5f",
      x"7cdd366eb7f4e7b3bcb18549f13a7841",
      x"94eb12aa40dfe2b7617817727c23658a",
      x"619158f762920e40ee4e2117e1184523",
      x"1031a6eccb0b25f536bf7d093ed0663f",
      x"430b9c4f28d8ff9bae3a3c9ef2883884",
      x"dab8cc10542c6e4880b22d1e220cf408",
      x"4d92a93ec09b6b1956f1732a9284be0a",
      x"c6b0ad1b1f73cce74e917849511de137",
      x"0fbe2b35afc4b72ef387bf91a6f6ffb9",
      x"8740ceeb776e9f5f8f2cc66ad1b8710d",
      x"b0f39cac05262ab009b69b2922d5c2f1",
      x"183402fe8677f196af4ad3300b1e0552",
      x"be4bd275776e3341cca69f859ad809bd",
      x"2ada6eddefe3d25434310b8941ace28f",
      x"b60f101799a09d0d6f85a40097786078",
      x"8f0d881d023d8590c66b9d316de15f79",
      x"1162e27d810e146bb6d72c48d0e3a3b7",
      x"e2aef8011171c3b298228a3e114fa651",
      x"207041865bcdbce967efd674d0c8c3bb",
      x"f9fb6f4aaac7a700a077a15e9e70dda5",
      x"c6ed57c81d6be331745b47cb5f72b662",
      x"20c69b0af8ffcd3eabe6cef39057f4f3",
      x"d7816b60f4ed5b7f0543abf042dd15eb",
      x"72d60003fa00022065853fc2778ea1fc",
      x"c59300d2b4e9ad2732fb1a4498b26103",
      x"20a8f09e343531a2b6f216581eaed49f",
      x"fe1155273221c837c34feee1c238f229",
      x"02b55a97b7b374ed92a08a29f5e5f7fd",
      x"526512753cb8a81d56f4cbb8d280bf61",
      x"fa0655c8babbfd9e9a5e6a2f6f9af0b9",
      x"66daff2fbfd5da590bce366c5828a246",
      x"08c8a819e4bda0b0094c68d3b7920286",
      x"e7d8ce949ddc67847e8de3b99deb330e",
      x"d01b618eaf07b72d3106eed237b3f30b",
      x"13c4007a402d457b169b00882444b3a5",
      x"4ed2c5d3c37156a490ee332b7953c86f",
      x"198c78086a8eb5aa5afb0ff6f10c70a5",
      x"7036f1f208f0e769f861420cf3cec178",
      x"20428c9446084035ac82c1ea1a6468d0",
      x"00ff1e0bd1df00b1bffb49a8d85eac0f",
      x"8860bea550cec3af95c618feb3f77a9d",
      x"00399dd8a2e9186145fd93932a9c8a0e",
      x"c9c63bd66339b59257b8c6d67ff94bea",
      x"ac421cae8ded300a3b3d7bddd880ba36",
      x"a515cbed068645f06c91f51819c727ac",
      x"c0c7995b7586e3493e92718513f7c49b",
      x"29bcec906692bfece93ef60054e64514",
      x"477605106318f533d8309b9aacbeb62d",
      x"66c7242501c92950c4dc64deebea0ebf",
      x"d2085b08df8a8f590e876159b45a7954",
      x"f65919c9673f2cdecdbec484635b21e5",
      x"edcae0558ede68ff37758f63ab60d66f",
      x"aef52681449f950d8729f7b21c063807",
      x"ac4b7951bda4a55a27e471ff4dd52671",
      x"9677f37f23e569e9cc006308fe490c59",
      x"85f0a20d5e5e967b9a388dc13a2be69a",
      x"4f70aa1d7d9978d952f060b1bdd73993",
      x"7d06ae233019c829d8f5fbf2b2d0f385",
      x"0a333616cede4bf33f74b4b7e988a8c5",
      x"6e6cdef57603597d0ae47724695cd464",
      x"81e049f23a14679b3662245aba40aead",
      x"be3a4130f14bb9f7fde883c5d027ccd0",
      x"4f07da2d497fcd82ced65aca0b9d2eb8",
      x"2171270cd26bbc7d3319a3b2d2af7431",
      x"bb1534e8fc0cc9be272e9c1ebcf4d471",
      x"722204a5920bb761d6363d8d4f1a88f4",
      x"55f44395c485bb218d1d5a4dcf7537dd",
      x"3e8f68a1d1a9caafe5b7ee65785b9cd9",
      x"add7d51439b822ecbebf31a9b261e00a",
      x"0e0c0363ad599eed17ecad3b1625532d",
      x"89d7778541a76930ed5ab8e997ee274b",
      x"4aff93ec988bec653ff403e75d0374d1",
      x"8df7089e11440884fd405f978f7de556",
      x"c1bb4060a5b5a0b9156bda092a8dd643",
      x"d4ac7339890085b1cb91f570463549e9",
      x"009c583840032708bf1c2f4f1f1b0df7",
      x"e85261efcb5b70be8fd61cb5acc718c6",
      x"2c16e352f83fc0f2d461374167ec7750",
      x"79fa54af4e44575fff6e5d18988326ff",
      x"8b9d422a236910b0c310fc27407db34a",
      x"bcc38b2ce0cdb8e5430b211f637e2234",
      x"3423811ae4ca05a0c4ba149b33630aee",
      x"cc542d09e0cc725ad7fb5eb4a7204ce2",
      x"feb789e2aa0b00bd2502b32124220dc1",
      x"bdc1b7be3d09b59a9d29458176ddd210",
      x"ca01b0730c8f4c62a87539ec21b5876d",
      x"9148d36450e073eac57f65cdb71a4822",
      x"690ea9f804dfc866323bc1d80322c21b",
      x"15fc85c53fd2e7697856f18cd0a04d28",
      x"8cbe35ff9fb64f2d26a3f65fb6da3069",
      x"213f0361332d3e8b6f7adcbdd917c1e9",
      x"dc203c894dfb652c89f38392e2d84da6",
      x"a6b4bb555f99cb88b872c2c1c8a0d420",
      x"78ef3101e9f88283984d814e43cadd9e",
      x"d1ec6e79b993c0bce6fc2b221da3ff5c",
      x"53111255cc411804b3cc929720e47946",
      x"6fa7f78b5b6633ebf857761fa2d886e0",
      x"990d5fbe05ee649fe75d3a51cf4cd16d",
      x"718a91984a4ab2ccbd1aa6c4606ed2db",
      x"1aa139b5559ecaf9fc115bf0060848a4",
      x"060330e43a1f0ad1d72cfc5f51e30d5b",
      x"92b325ce30a9c1ec57846b42da1f6398",
      x"3572db72aacf6c51f01332614ec84d9b",
      x"cb319be534ecac7f2f65cfff10cc6835",
      x"4a1113631ba6675df8e37d04b37f3a1f",
      x"adc3183e4aac84cfddce5802102e69be",
      x"1bf3f9dfe6e5a299b0b3c04916ba32c2"
    ),
    (
      x"9cd662564dedf16128a018cccde39b97",
      x"91784ce8da112eb19d7da390112ec52e",
      x"16ed8f8d75a6ddf205715fcde048b4f5",
      x"def71c2ba0d96364a8c017adbb7e6b62",
      x"f82217770dfffbaaa9ea6e0bedf57572",
      x"63aaaf7b9d7ed2ac1017b0751a83fd76",
      x"6e3425b8bebf6002411a25eb04a135e4",
      x"02d0c3429b199b687c155fd8c861ed00",
      x"e4670eee5837af794028f4e36b724c72",
      x"e53991ae6bb169c7dff604fe5d05fc88",
      x"fd655a12cd8b6935c07c57fc56fc87ea",
      x"92eaf36ef2bf9426fd67518469ea21c9",
      x"66bec1b6854936f2632e3762e2602d87",
      x"6de9f36fc0220477166976983b7de5cd",
      x"344e016dd586c57db745823156f01ad4",
      x"f2336426e2e27cf67c2b3d9ccbc7fe42",
      x"8124007110c6941c050adf4367e0eb4b",
      x"eabf44d4fc6cc02342f95ee921b7c1dd",
      x"0afc0a7499250aace323b9912fe26051",
      x"ff18c6efc3f66be33c923778ddf022fe",
      x"622e08be970786a782ccb8d17c1eae2d",
      x"3cc4c930eb96142f918d8c618b6f2e2a",
      x"3cfbbeadd26cbe1f7a3082922ea36fb3",
      x"d912894c56d9b2e2d30e8932bebfb820",
      x"c207cfcc7df1032d71a611569f33795d",
      x"7c8744d38d5c95e477be08436a366cce",
      x"f6d80bbbc4a2bb906f131c3868e97e13",
      x"b57bf796aa93a75a1b9a44709c04b991",
      x"665abf1d6883a232502ec147fd83df31",
      x"e4fa1c7686aaeb554357014553f08c6e",
      x"a23a0c6f33a237c9327280cb8afb42f3",
      x"4602c2e026962db8e53bc0e36e5c2e53",
      x"56f3694bf0f4e4c50eb262842e2a2dcc",
      x"f2bdf0d68d4be12d4bf8fc0991c443cc",
      x"8f2a85919902aad1734296e852128738",
      x"fa85d8908e742e108f54989ffdb67b36",
      x"f089a641f8f2475a40255e4de7ba273d",
      x"d511918ca896817caca7d025043398bd",
      x"f8fd257a397e66032b4763e64ad9a6c1",
      x"35166b89d303a4b8eaeca5822a0360ff",
      x"880d0aa7fafbd79d0ad24017cbad4ebb",
      x"26cc4a32ed591ab88674c33654aba398",
      x"263790117eb3fbf5f21013877e37a8d8",
      x"d1e0cbb176e3bda39f7d2548a5fb834e",
      x"570a9356d41c4fd2ba356d702f80dea0",
      x"8e99e9dccb4135ce95bb5d5a42ef9557",
      x"8c224164ac89d9a23bcd3a3506ff2536",
      x"9d831f709d014360e4a0726877b64470",
      x"58b405f142872cd426bdeda7e1aa5a20",
      x"b846ebb31e73a309ccc5230bc5e73d7b",
      x"5a691fbde8e1999f67cec25e27a26464",
      x"c6707407988392fc9631f8d91d324bae",
      x"7f0bb068b8eade0f01c8a2bb326f4758",
      x"2bff950cb85a2ff263f80d228e58e646",
      x"695d01dfd23eb6a09d7369849a055a31",
      x"3544e6db55f0a84c8cc99dcfccba3397",
      x"5972b18abe389c0c0fe649eb5ecdfe81",
      x"94ca612602167305d81ab90a11253967",
      x"777e1365dc202ff152c3d149b1286721",
      x"78878aee75819cff41ccafec56044381",
      x"feea3c2517616eefdfc8ef8fd23b8521",
      x"3349286e249fdad337945aa13fa9f6f9",
      x"c4da168cfde8f58f05e32ca6c4d40488",
      x"c44181789fd6788737b3ff8ef256c6e9",
      x"ee63f1d5623597ad334e02a5c97e4ce8",
      x"faf2a5901b50d36fd4b8a0c859d584a3",
      x"36a6d5dd20b3b799511cea1998badc28",
      x"c2aad8225f5bf43ae0ee54cf93e4759b",
      x"ba435e3b9e16dffc94f449b7156eae54",
      x"7086af8c1579023c9297597bd15754db",
      x"70696ef0d2e4efb4b5bfff5d79ce7e81",
      x"359270071042c9818cf7f5f69aa2b8df",
      x"81954b390434d27f3fe1eb3d74dbe631",
      x"ed0685f77fb1f404052637923f8bf48d",
      x"0e3dbcf592d21b4ed8492cf82fc307c8",
      x"de47687ebac4112530d05854dc730d66",
      x"edc2eb1af17c647fbce140b70baa169f",
      x"aaa4161328714a64d539cae66d690481",
      x"7f6b44c3e6453af2487bb7033a7a0cc1",
      x"a5f5c5d7e827e3017a4ea7fa8c92589a",
      x"ec6a3dac71e9bd0d7bfecbaceac43cfb",
      x"5b1a1f782de2514a8209165e55125fcf",
      x"ac3aa9675308df69e1027fda316eaae8",
      x"b62998daeff1bce38faf9eeae0883c8f",
      x"9edd19949e76c1fb1dfa1fe636fd564b",
      x"a755ce17da24032e72c60e5a69bf25c7",
      x"51b25bd57feeb65fbecae7eaa8628fd3",
      x"b3654bb7a984d11b0b71e3fdd71b4b25",
      x"cb54b12ef2518a62f8a95cbd11734e60",
      x"42f4f74eda1da8de6e98808e9ac78bf5",
      x"3ff3c723064daa5e5c50a3a82565173f",
      x"1de18f658de948a4d22ee9a29a76c848",
      x"af621a97490d6682279ec5b08bd21151",
      x"a7f3f50d33d5e9dd4333c25c1189f319",
      x"0e83a639be5c6628f6605749b762628b",
      x"ae3ad23c6f43a8c3548ad441fc471502",
      x"7fec2392ccac543582c0b28c562a3581",
      x"2efbbfecd3a2953244b896d9b1a1e038",
      x"58fc3107f64ff06076be1202895a28f8",
      x"d7a41751861f7e3e56c1c8e0a1a58528",
      x"82ef7ef9c8074cf565ea6b7e316a7114",
      x"08edc75b513b7b0da62a4450f15d1cee",
      x"e4a300e192a525fc049179f92ea80ab7",
      x"a37b50a50ebacae9fcc392b7b180b40e",
      x"b905804f0c92094efc7d80229ec36708",
      x"0bc4b6c08fbc74ae1e82cfe022100eaf",
      x"13c5d7acb0df664defd0768b8c1da136",
      x"4635faf6147348749b84f0b9565bf993",
      x"30e3142fd49c52cc69edb683b9562750",
      x"b2bc420c21357df8e3ded9a34c66a8a0",
      x"5aa19bd77cb6b2b5de191c72b3625237",
      x"a875794ff70b04d401505586221d7bb1",
      x"5c2c5ecad284ca94cbb290d5a902fc31",
      x"290680ca25dd64d74be9680f9b026642",
      x"5ed42460a43a2aeb6e06fe6700c2d7eb",
      x"19de7cf141d96240ab542e8f203b45dd",
      x"cc60f5453bd25bd332c31a1a3da3ebd2",
      x"b5d156a28ecdaf830a4bfa956dd65708",
      x"70d77cdc01ec0c09b4a57ebd2ad2a198",
      x"0d4aad7286dcb8fdd743aa9516c8527b",
      x"c03c65317a34af305764dc2261ee129d",
      x"0f45c22eb63ed4f6c705a12666385955",
      x"65b1f37c37d9d4c8c13de734de2b2253",
      x"68d86c9a09af9eb7d47b07f0351251a9",
      x"52b188eb4f51ad0e30b6fe2385058611",
      x"e40e1fbca8e7511756a901b33f31c1bc",
      x"85c9d5bdbdf6b5f608c910b244f96000",
      x"5101e09bada9a0f41ae79ba396073458"
    ),
    (
      x"6fecb12879a7d00b970fd553ad5b1e90",
      x"27b6cb93b6f860a4a74e3101480f15f2",
      x"e7c5eebff96df1abcf0c746fcc56a375",
      x"b0686cd11cc1b95bf6b6c5f2c98ed60b",
      x"79a35f2314090b0b2364d98b2fcc7ca9",
      x"578333ec70896449ec42be9e1f0126b1",
      x"f21441587738835b867e98f6d3d91059",
      x"21d763cf86d3803a1765501537f0ee1c",
      x"9970aa41aaa6a4b840032aaa4f4745e8",
      x"622d404887b87ec4192a18899efa22c4",
      x"9468c76c632fa2235c3c84ce685ee302",
      x"b335a000ff2f3e77957346a20f9381bd",
      x"556e31029649e4fb9a5593f2965c011d",
      x"cdf67d4376aadcd5ece17d2b8ff57b03",
      x"d6188204ea68ff51682ec1ede938d4df",
      x"7a2a02f35917f0803902f07b3180f377",
      x"4ad59e2126a4c636d7cdac9b542d5ba9",
      x"8c36622a016934a8ecf980b717d910f1",
      x"973f115864707b34cd4d82e9be81d70e",
      x"b53980c162e873cc1523a3d2f91871aa",
      x"07e1d3dde868d14fd7a65170aca6e2e1",
      x"7fc8da14807ea689ed5bd980fadeb20a",
      x"4656dd5bd6c221a43d6c3fd3ec3216f1",
      x"4581c5e6c2adfb0e63b80f612a93b9c6",
      x"3989bcf4a01706e9415d96517e16bcd8",
      x"c0fc32aee6d16e62d5e0455546d5a4d2",
      x"f5e35dc40d5a406d56638225b151c9ee",
      x"2e50f89c0f9139435b60a7f1cd8d7138",
      x"c0372c9d7ecde7a541638309ffe1afe3",
      x"386a534be1df43578b938db0e9bae9ff",
      x"bf4b447fdd0bb6041c17132fb4bdf22b",
      x"d7c35f3c6686d0f82298e9607e8cc8a6",
      x"5c426c5ef2cf96209d5931291f60ae72",
      x"96a31bc881c8c6c315a7e1dfd79c577e",
      x"ce9827d0ba00952b4995487d78b98ca9",
      x"1bb54540bc563ac3ddf1c1722f3e7d47",
      x"547eafd76f14cb6de223b5d9033f406c",
      x"b5b5f2d90eea42e79924c4b237d4986e",
      x"f1b5b6a8727615ecf016b8118309c937",
      x"16083d00ea5a65f317a694e6ccfeb3f2",
      x"2de26b6902e0187fe66453510911fd6c",
      x"843de9ab7c7431cd9ee53d2795d593aa",
      x"7387a8310ff9f3d9e83d21a26ce90331",
      x"1be5865c95fffe5aab5cc427d24dfcca",
      x"fe02157cfa939f6aa869a4a7c658d000",
      x"ec8509fd3bd6bf8c771e3a3c8e328bbd",
      x"d76aac9f1bcf1b8c2d15a1cf44c45fdb",
      x"a9051a688c0ce0cfd99b3f317031fd63",
      x"79f4a7ef67b08fc8ee0871c7d30a96d7",
      x"958c94865258bfe4e26561743f82e6ca",
      x"1d7cdf476f5f27446e1acc0e0e09d96e",
      x"9029e62fefadf4351f948bb75989c78b",
      x"153901b061ac88ea5593e2fc7796df61",
      x"ae3950e9e6fe7ec0b8627476ecbf26d6",
      x"256dc142927cecd5629ed07f5312eaad",
      x"30f74587de63851cb6eafe0be0ec1069",
      x"01605339dcbb90e0cb1e86f913e3aeea",
      x"f2ce58363b2ea08f154014856743b226",
      x"8c915aa9012f68c92ef31f264675f9a6",
      x"fb45d9e329e4195032f45a19e27451e2",
      x"e1a25e999b9093b3c183b07bc668ddae",
      x"48eb7c8c7046d039e70f7c8076590294",
      x"b07aa54b75dda3bf8ebef5bf87ce41fc",
      x"7711ee097f3c845e1d1d05c978a9675a",
      x"4b8b29f3289ccd667916307e6e911c55",
      x"c30024cf7d1e8bbed4257de0b9533e85",
      x"5b975c6048f9fcc059a0ba88d3a1b426",
      x"cd8dca30dd13d1c6c8d0250abef50145",
      x"4d79f385c2b818d36963edb21eaf436d",
      x"1bc362c0b5b746795f4c2d4ac7204213",
      x"90595fbc2138f1e6c5542f1888e2269a",
      x"88f3fa36fe771180a6334ce6d7d016a5",
      x"88490177f75c5b5d4e18af5f3e37b91a",
      x"3d72cb0bb113a14f22e32c3ac2964c51",
      x"7693b65d884b479ee809afb641d53887",
      x"90f269da40f113dd75da5e30a956bf0f",
      x"b4e6aa3571685be39ddffce48dcd0fb3",
      x"0fa392872498591f488220c7a35c795f",
      x"6d3b0eaba75a78ff63019f5f126bd554",
      x"c0f05b1f0d638bace248651efd437819",
      x"b1dd3c8c5a9b9682d49fa486e56aff9f",
      x"93910869ceff9ce355cf9bcdb84d0030",
      x"2fd9c4f2e9095318bcab1953a7852491",
      x"3b645cfa62ac5ea7e04afbc1d605f83f",
      x"7d2dde0545329405886cfad1f960d407",
      x"a718a0076522c0d74c1514f3b2eec1b1",
      x"14500fd02fa2e00a8548d6e5273bc335",
      x"b219340bb687f3e3452c6b3f26e65997",
      x"fe78e7e6275e57fbf31a904720b1fde7",
      x"b9dda5477bded037b90a524ce92f30f2",
      x"4a867766fcd8ebb3012b37974f16a634",
      x"65111cb0c988d0a6727be1e17f85f503",
      x"35de56e7f12798493c95910f528bf7bc",
      x"967403b8bac1e9b8cab92a8c57731412",
      x"45d912072201689e84988f6433a8318f",
      x"1d2eb4243d3b93b16bf45db400a14caf",
      x"22bb6e9b7298db03e7e522c1960559dd",
      x"f4fcfefe9a360805a6eec60b7034b992",
      x"a3872b90d6c0a20914db6182f1220ddc",
      x"d986b4765b0fcbd809b42bf4132df6b3",
      x"a0468ef73d1fa7fefb2da99472284d39",
      x"268c7700557c1cbc9f56ec2c697cb27b",
      x"84290d426dda2fab7304708fc5174b05",
      x"c7799cb6d6ab86e41d8e5e171f2e3816",
      x"308f6df7d395817824e11e290fbd4211",
      x"c0a0d8ccaf6fd598292cfaf92b0ab0e2",
      x"8a878a0e3583554da434be5d085ce23e",
      x"957a58b134eeb458388b6770bacf4cf2",
      x"e885a5b95f2813bdbbb8300d995c2b5d",
      x"02e1908237c458a692ae37abf5e25c0b",
      x"77566ad4a28ca43e795e2fc713c420be",
      x"eb521dd5ebe3bb2d69149ad2e44726d3",
      x"f1d60269d1daa3ac8436f8cc823658bc",
      x"6beb6b0fb2922cf68e139773ce31eb69",
      x"50b60b3480d3da7da02c5875683ba674",
      x"f55daf2395b4bde7b5b1f8f7947ed141",
      x"80083c2c75a354a92a29089d7194606a",
      x"61b07bf2b0cde7cd169aaf869b509506",
      x"dfe6621671eabc2265e5633837c8ad20",
      x"d27f78ffd8b4ab9da2b70ecae4b4ccaf",
      x"e69f22f9ebfd2015f5a93bef6095ff1f",
      x"352de037d25a3c1214940024736ab878",
      x"5d6670b51a166485685bd51c1bac89a2",
      x"91ebe4a02f64ea3f4a3588b6b7836e7f",
      x"e0291499107ed1c7e67e612448190a65",
      x"5f3617927ef0219bd74b353d00f96c8f",
      x"b7e9ec0cdb2d48217911811de9e72ac2",
      x"cd6d900d4debbcc6ef4528ce4c87e1ff"
    ),
    (
      x"a578bc2a13dc40e9486e1a9aa92e7498",
      x"10ab610f48aa15bf361829f67d879bf7",
      x"472021743592e95dda58bb46166ce618",
      x"593628d063f101d6102198e8e547aaf3",
      x"add614940dd92fbae43010029e775f89",
      x"7d9f992670f63465e0b9125876075986",
      x"8aceb851360667fe3a585ff7690e3a09",
      x"829f47a93334b7089bfae5d58682bb69",
      x"0598fc885349a625a03948b62e3e4678",
      x"a0c57ec8ae010a0ead3e2243f5ef37df",
      x"4f695e0ff2f7c193c353c74969b767da",
      x"ec1f9e6ad61751b00f3c11b1e9af7daf",
      x"1dec62dc181bb4d17f4a06c4f9c3a968",
      x"330f427785686ea2135448909ecbadcb",
      x"41305926ad3b519d5a9eacef0367c206",
      x"6f17d585147adeb3dc0c56f0343c5d5e",
      x"46f9e496710dd35fad2884eab144eee3",
      x"9ff34914084e9f415e2960d62f06b03c",
      x"5aee5ef05146532750e0aca2fedc33b0",
      x"d1b158657a9da8b02f1938254de6f4b3",
      x"f6971ee74715812d9591fcc232ec1dab",
      x"7f959605da7bee8141cbe53269cd3f38",
      x"a6b29631075a5b485a542a7b024de589",
      x"b527a181a91ac4da5c615098e4b188c5",
      x"8fdc55b131a9aa2b482c34836241fcea",
      x"2078ce89f40515636d57cc72977aa2f3",
      x"22a1a3e4ad3cd0733d2e6ff538cbe5ad",
      x"227e4e8d809fa14319384e8daf1052ca",
      x"d30660fdd49992231d015dc8714262a4",
      x"a7b48af38bcec257fb7fdd90bf652664",
      x"ec94db88fb1070f76847396a2c1930c2",
      x"1f368a5147d9400fce0ea863dc76eca0",
      x"328cec7625fdbaf35d0a20043851da9a",
      x"d5dcf2267d95334de5e6ad326cb77ce5",
      x"de3e44edfbddb0f4929c7aacb5c6d51b",
      x"55ec9e6f58a523d3582d07d721129908",
      x"f384012994eaa10f8a900b2398e29105",
      x"5e090cce0f81dedba981375a9036d8a0",
      x"afa5d9be1b498953816c75158d4a89a9",
      x"c099c517254d43cb8710476ed4758909",
      x"e62ef51cbf1709053de1753e712e736c",
      x"3ee1a3ede366bc96c8df0028860776d6",
      x"b9b094bf37389073a1dc7474b4d23a34",
      x"b82aec9257313d7ccb55f226b624f72a",
      x"4297c50677d6953d04bf3978a7108a44",
      x"1e9696f8821465cacd5d29e90c3fc38f",
      x"81db8c6b67ae3c4b8f1c24ede08da881",
      x"4be925064d7d30336aafe029614d8265",
      x"fba26eba726ef97b811235cc89ea2e7d",
      x"d053e5ab52eafb600fb1cd6f5603ab01",
      x"cbe000829631732fe6e81c1f4099dbbc",
      x"4d8a51b45fda54e2a4d202d1d58588ae",
      x"7e41c4ed31bf52fd20f3face77ff4a3c",
      x"61b363c63fff9cc743ccb08bafc438ab",
      x"ff9baf350202efe3b80b225910e560b9",
      x"4bfb1cc46c41cfdfa9aa13f0fd755619",
      x"999705ffbced65df12419e6e21bb0bc9",
      x"4fede9660563abfcfd0d51900fab9041",
      x"1714975bb12d1574bd646dded47501c6",
      x"ae2fe46d0734bc7c6c3e00073bb64c4a",
      x"d7d024af3cb3685859ba2a6f149f18a9",
      x"a0df04fedacde5526311b16f5267eb17",
      x"750638684afc0b1324445c317051db14",
      x"083fff97c0f1db0600db2bd1420d4add",
      x"9a35fc29d5628b31e2ee79b55a6dcdc0",
      x"44b6eff1add03dd42068173c1291afd3",
      x"0b08e62d4adcbdb5dd8a2c1449f27b5b",
      x"4afa7137f32fe1d07ccefa77a9222e23",
      x"92503ee55af032cef557f41a3bdc0be2",
      x"3075649f8fbf1531ecc56c2d19f0b4de",
      x"a35c8895bb7123a0f924ceb1c86c8e58",
      x"98a67872938cb4f9713976afc0574077",
      x"771e1fb3102d2e66ec704527aea9921d",
      x"5b2debf5bdd9659c80c910b30f9ca660",
      x"fb907d804ff392fb921f2699252cb8a1",
      x"b59ad77997c24df983ae6c597aa0d119",
      x"6263b3dee3d0323f222ab8fb15a5f1ee",
      x"fd31be79c75576bfce441bfbec59aa13",
      x"648500f81d7683d03a1be6e03d22f864",
      x"d9d32f9d59ae9fb4fb5384dcbe4c2465",
      x"076de08f07e9f632329f5bac773fc5a6",
      x"cabdb1d464c0a740ad0326a726629521",
      x"986eeeddcce4a54a448d3451feb64187",
      x"5aae7c25a21ddbb539460778662433c2",
      x"d5db86a55f08f9bd0b7eaf2ef61c373c",
      x"fb478b4fdaef78821fb69d8492edb76d",
      x"a4f19016498f7d9a8b4737c2361ff04b",
      x"2928bb280a1f858cd5e99d2032e082cc",
      x"61287e767a126096755a5f2cf1f3427b",
      x"e35abc24b07cb5ae0db0a1d2f373bf74",
      x"e094a7379ea8543d85bd278d29857465",
      x"99848ddf36113aaf229972532ab6d0f1",
      x"f0a440974efecdac76b08a2732b4a829",
      x"9f5e2e18c7fcdfbe87679a02be3ef970",
      x"23792cfd9436f46ef2e05816f511d28f",
      x"b7f1b8f8c5320599c9c4887e791be32d",
      x"8e5a5167fe9ae8589a94b63b532d4a7a",
      x"1fee498a92e2edee43edc571607506b7",
      x"6c8b9dc3fd453ed42bb6f34ad56ee213",
      x"9efa17f644710d6da8febf341c0bc3dd",
      x"2bae1ab0d17fad795308a7c26dc5fe56",
      x"f897dade576fde2d93753f36729a7951",
      x"5f741e6c3859eceb081f0f20a03882c4",
      x"68fa3ab8da0a7160ef7ae2e56c990a86",
      x"0f71ea9adf259f633ef7dc36264cf88e",
      x"2de581293d6cc5c8260ded1e84e9b89a",
      x"afbd53d9ebdbc8112d17260cb55df1ef",
      x"c3c5a6ef422120c3ae2a414ed346a7ee",
      x"f045d31861b20484a82e717ce87e3f26",
      x"234bdb9fe05438f47670139bac93095f",
      x"c0bd1f26640ac449e8486a607ba43ae6",
      x"a7c9bfe7afe649de86decbf822ae4362",
      x"835d902ee1b5591d503823266ffe7e1b",
      x"696bc7ebbef46b8d4df7038243b4bf01",
      x"c56f03b8ded4f45f510c15cfc9d1edd8",
      x"556f49d24cb17a7210f060e61cbfd1af",
      x"2c5adbd7cbc24b98268420aab865ee03",
      x"4abe17155c5c145f5f041099b4464b49",
      x"d55af7e828c8ec963d09a639c49f4afa",
      x"67d2c517b862f3cb28cffafcaf965163",
      x"bd376e97af2d74fb8d346e810988f80d",
      x"de66887347657d1c0f314d8f34daa575",
      x"9a5dc3d81afdcc5d0eb236bb4fec49ec",
      x"f38ccaf56858d0e22e826a8d9dc58dd2",
      x"27eee3bfa2fef7fe0d88acb749f7be7c",
      x"e983f71ab46cee00150f9c4328fa24ab",
      x"80d7a07a3b9fa7aba1b1a069e961263d",
      x"6c59c74b20bdd5064149b734b2ad2b65"
    )
  );

end lowmc_pkg;
