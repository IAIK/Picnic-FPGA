library ieee;
use ieee.std_logic_1164.all;

library work;

package lowmc_pkg is
  constant N : integer := 256;
  constant K : integer := 256;
  constant M : integer := 10;
  constant R : integer := 38;
  constant S : integer := 30;

  type T_NK_MATRIX is array(0 to N - 1) of std_logic_vector(K - 1 downto 0);
  type T_NN_MATRIX is array(0 to N - 1) of std_logic_vector(N - 1 downto 0);
  type T_SK_MATRIX is array(0 to S - 1) of std_logic_vector(K - 1 downto 0);
  type T_SN_MATRIX is array(0 to S - 1) of std_logic_vector(N - 1 downto 0);
  type T_NSS_MATRIX is array(0 to (N - S) - 1) of std_logic_vector(S - 1 downto 0);
  type T_RS_MATRIX is array(0 to R - 1) of std_logic_vector(S - 1 downto 0);

  type T_KMATRIX is array (0 to R - 1) of T_SK_MATRIX;
  type T_ZMATRIX is array (0 to R - 2) of T_SN_MATRIX;
  type T_RMATRIX is array (0 to R - 2) of T_NSS_MATRIX;

  constant K0 : T_NK_MATRIX := (
      x"c24f16269830180b15c295c21894889c5a4993bb70b1c39f0237d95c1e832002",
      x"f640e924b648d06edea78046da1e78a26d71fa9440860faa4cbc257c47d3c096",
      x"3d3695b840d6075fceb9a455d71b25de18836fcc47d605fb1fac80409daf26e2",
      x"8a271257d44205a985ded37c470836d74ad0e971324e3b862a3963a5b9c4f7a2",
      x"df2eb407ce27572ae41fdcf686bc11d061599c6db147d4e978eb04804e15ac95",
      x"b0e074126637510f3107c01c2c656372546dabdd57d3cdded8de215d348956e1",
      x"77cc10270234b8eab976eb6a7bc14c9e73a12c6b146c71f3aac76cd76f8df8c0",
      x"7bbe18d775183d8345ab2f90bc3dd0febc5bdd2860af20aa44ac6b22d5c5e32a",
      x"830d1ab541a7d07a3d98adf8bc3e15b30a9eb112e2ed341593fa95cc8f83a049",
      x"5d25139cdae197e627e4d26db6d50ae2294a8e9ce384d6e3f20965fb2edcce00",
      x"7238e686f74aa3d30d735a6e88d501686e8a54c7583996b20e7115685cb51cbd",
      x"5ddd8ba2053277a1c6360cf4db4378c956836e9514d0d9c3451432a14df86dc7",
      x"3a2d05e8546d93c5e3ce20a26c95dfab010a1abe69d22566badbeda186132eff",
      x"2b0ce15778fb6c90ad140434ce367aead4c659e347822d26275dc92cc3a616ae",
      x"423824b58072d20426cc26bec22f1f3a5465454a7e864bdbe19261b5c27e5cb6",
      x"db065668b86a73d41197250e1f667ad3447db4b113525e0375cfdfc9471b94e2",
      x"f9531a29cee0291d83b2cfbee6e9306e099ecd3146796c28bd8cd97803eb156e",
      x"a34178670211bf883a60223864b86dd9294a14840a9ab08a3ac4a1f44847bc55",
      x"38a8892657bb861c65257754b87b9d297b41b2db0d8ed147cf7e8a958e5ecbf9",
      x"25495e9beb966e72e83880922fb678c2ff91e581b563f9f2b16516321e12a707",
      x"584c3e22cbee4b51cfcfa8902c657904f1b0f6e9f37ec763f890e30e3f238d4a",
      x"8e5b76495103200a6c606607fd4842ebf5f2c826474028e9af9b169ef27cf5f2",
      x"45c2b9cab066791dc533a34ec635f438f7627c146e04430918ee12333ce27718",
      x"dd6d8a359b033f33053da7878b7ae6bf0d340ca47bd549c94313f318ef671179",
      x"1886654059c80e73cdbd9477835c0f9a069b6a323fce5ed7a771d981f4080073",
      x"ac58c02e866ebc9abb0af12c99a746bf35a0b342bb5648679cb4076055c83fb8",
      x"4812a840b13151f53d93641d7c300fd1219be4b8cee9a5fb115fc08f623cd847",
      x"15de9bf62f74f7844f39b049712a8f88d7064f2c8cf6f4252b4b31564e352705",
      x"697b604cc8678b12f3394e0ec80120e2efb8242270ab8ea7c2af2ba5046add11",
      x"42b1ef0166f22fb094bdc91abd6b6a1bb56aaaf6d440ffade3dd959ff43c6139",
      x"2f7b1dc3d1f522b03b1bba8d093cd4634459162ca9d1b571feb93419fb3ee9ff",
      x"9c60f72528fedcba9213efa8eab9c3f9427ead5bb95afeaf50aefca690790061",
      x"00996f849641a73e29292a1cb01d0e9426cd1ec0167a4bd1e93348f0deb0bf19",
      x"499b674e47658d70a9ef34bcc5eff568c4518440ef0c38dd1044bf14bf529b58",
      x"3a261a45f9a2629ed52f5c5060c2ae87a7929ee4bd8cc177b0d78f7d50e159af",
      x"240edfddaa2cea8e4466ce493fccff26b3a60c883e7a3896becb9df8e77584e3",
      x"4404dc19db5f5650f18fd0f2164e899c27a7acea565184aef342742025c05df6",
      x"a460f29d89f60a5bbfee3ddfd1b6e62bea592421d0a14c5418b1ef9e0483e777",
      x"09c1fe7d3c232251481d0762aed68c9d9d2125a96564b258c6e087289c9e533c",
      x"7eb54d97df60a20ec4efe0f90c2e482610063630efdb6538a965f6603598b223",
      x"a7e14f3e7eb11b403e3d91d4d5c3fcf66282a4861d628ecf089e942b09954e17",
      x"d5a6234032fecc09da57f7c288a0ff2beeb267dfbb6869b21a757771d71eda7b",
      x"261ba5c44ec3ea425391146e389041b221dc68a2ae13eb1124ef34a18c3bd9f9",
      x"5aa5ba5ce9fb227c597e4ed12f13439a66ffaa10876d90967083e6f3d77dfb35",
      x"f1702c44ba077301d88a8a30776e2d4b26bd61a6588343c936cc0b6a116ab01e",
      x"dbadcc7268a212e12a46fee16d4abd86e08fb1265634edb47d7ff6b9597c80d0",
      x"01b9615abf0c900b78ee086c8247ac98f70227697e50463e085b5c8117efd76b",
      x"5672aa4ba762631a073850d035f03c7958d7de79f716d00edfedc4bad6d83d8e",
      x"e2eb32a1779adbb71ab641c076b3699f2c672237cbd5e673ab97346eceedb5ca",
      x"ea77abddb3ab8d1b79226840ea7ffafa4a2a12a2bed46affd8d3ed5383d37cb4",
      x"aae004edcaeff2df5a4d5f7537a89f7f0c6393a7a3f4056e9f71a869d47b6da6",
      x"2f6a4a14d675af4f62a09bcddfdb7310fac2a45514263a9196ef2e1854eb0f78",
      x"354ed7d5f3c33d10c4037386ce9acd68029be252861c6a2e0b2299bbb83258ef",
      x"31dcb6b20f2731df54362af0ee3f8064e0f4da0bcadc1fbec7c6cbf539dd3894",
      x"2a76fd866e09fbc9802ce6753064b3086cc9aa7ce7d93b007f2fe87f95927906",
      x"57fe468d84b1c0a65029eec408111da95b33bf49c99a4ae8b8c7f27575194766",
      x"13d58147848e05bfba9f5fea9df07061dc50003ff6ea21423ccd4d87146a531a",
      x"810f93c83ce59864cace66afbe4cf9159198d84c55e458d2cbe42f6317b104e0",
      x"981346e4523967f263748511de88dc0c9b09a344f7c9a12569c61abec116cc55",
      x"fc5c2cb25e5539545f97190c85d0e66bcc431aaa731e7e46226736a500ebf79d",
      x"7cb624cc7abc85c94928e9b55c764936b208a64b8c242d82c509fbb8e2044bb9",
      x"b25e824f997116505ecaa3fd2f3bd9af81f463e9e013b897903810872a5fff17",
      x"904ef3b39d9cf163e470978508d8cacb6bd6ec395aec35f701ebb9a6c266d4bf",
      x"237985390713a7dabb4a1a33cf5ec359c5c2befa603b51ba818bcf1a00d2dc43",
      x"14392f4a50527346edbd3a666245d64619a5893e1c569d1f97293a1557d6e835",
      x"fd7ef5fb9d113f8c100f12d0ca596f8a916e16115fccf32b670c268dfa5ddea8",
      x"036a19bff4ac95b845d4812836899e1919acd429fdb38b0059673e4b33c8aa62",
      x"11a74e863851a986d32f334196d67819d34437eef1103b48c1a42116752e1f5e",
      x"f7117fcc9d5870136a939ce76c0886c5c315447808cdf6704ca90abeec77d6f7",
      x"dfe2b8fe2524c95a2444597b96bf3c304fb35d20d14d7288c5ac19d57e6e3809",
      x"4dc18c6aa69a90106a8de8827ecdd9783247ae8b6a68aeb56df09e4c57cb1713",
      x"2c3197916fdee6480393ddfdc9786756819099bc0f14f02c6080245e9c81ac8b",
      x"8fa1d9857a8b1c9a97c29f03af6c8e48be8c8e31f206b2a6bafe921af83bd522",
      x"40024e38234de27d7186edb79e0d15ee96050e0b4dbff8faeb3dd93def86b649",
      x"5f5ddbab5d343a445b111ff0aec77f137cae6003e97b16f39f22fa90267b56bb",
      x"d6a0a3bed34676abea4bfe3e575fbabe0d45141f50b2e2577c86a8c3377280fe",
      x"215bc47fbba2de00b78c0d6a655579fd08214a9b0bcf39040d1cc5cd25640a06",
      x"1d1d439947c5518111299d4cc45aed3d2850df28c5361f774e7fdc4550a312b7",
      x"687fdf52ad40235560450a0789abf5480c21f6fd5dc544664e302bff6db81592",
      x"d2a187ea1cfce06074d796ffb9ece0b71895009824cd9076bb752ce8c75a076a",
      x"8825007263782bfa7761e87bab61f5a4fa5532a4f464f2db6fc406d30c7fe15b",
      x"79a1105ff7cf0125f6c9b44165afea7572d6348a73697937d8c400a5985a6a54",
      x"86dd9a95675cb82a557c3806de4e048c218c2d43d1d6276ac462890d70c7dba6",
      x"2fdd71ba44fa4caba99ba6b4dc9794ccbbd0fa951a38c3465b8dc34115782072",
      x"41a6767be5fbafd83fc5f0bafbb4d7025b82875746bf9596aabc6a6e572cb39d",
      x"b406cd54971d48fda82b563b89ce6b50cfbb9ca77c7444946f452d9139b1b59e",
      x"d6ef21482156f6a2b361983bf26d41359288c03aab308fbf9a7a34aeb4407715",
      x"8986be8ee9b8f36adf3012aa2a619ecde57e9f1e11781ed3a1e2a1a3a9b1195b",
      x"b39d58f9fc03ae17e8c785dbf6555633f92d8fb932450c4cd7060568c003cfb7",
      x"f931c22e85f8a9a2a76fbd30d4f50adb0b9dddd2d8997716512dab8314277489",
      x"da3960fdc36656482786206945529d4be95f900aa1919a483cbdf9c7d0cf0ce9",
      x"b92c60e94886121c4b2d219bf904fae5ea06df7b793e5498ea8836aa8c743a9f",
      x"18051b67ec7a55f9587bf6f82685865c9bf847d60964351e255a79ba57e88fd7",
      x"c99d0eff7bc04f823e874d02eb475fc8cd98cdc520354c89b3bc206c91a1f4bf",
      x"95a2b0c6872c24418a01f2f05a76f0a7023064d492bef254f7194734c32d5dde",
      x"6a8977cc399eb408cdf6c9540079a9ee3f12151b43983fb3c9d382fdc27f2a27",
      x"c33fcef9c4fbe2c5902393a5eff6a8aa67e1111d9d7db4b3d4a64d02f8335762",
      x"c1776520ec7fc37142faea44c71cf248d1c74679db32dad31152400cd8f25de2",
      x"ed80fbbb08fc7e300933e609ba903fb8fad082c26b843002446344e0619b3175",
      x"6afcab88892f7b6eda5c25959c854194b20d0186f92b199bf29a574b308f23b4",
      x"1b02bbb0be7a9a9bc175c99b5b02020263bbea84937f5e91a597c5b1ece784b7",
      x"4e567d7b4524bef27ad261a20e81dff535ba83fa742931c9f726287b5615651b",
      x"0a60bfcdfd7430d1a4cb2908ef44a7feef1d0bdcb208c4c9a3f624910edc72a6",
      x"16472baf01170d8dfb16f57b45baaae5dab527117bceee32205b0217034985ef",
      x"cfb2e3b9c99512eb00e119adfdd771e6fc115a172ff564278f40186b51d5fd7e",
      x"1a8b06d4283d3ef90bb8f04afadbfdf2e4bbe44695ac0a53056abbbebf2d24c7",
      x"a513d6803f7a04e20571328d3b5ee408c82fc8ad591559beb69d9be896aa366c",
      x"cb97035fac89616207c8f233abc7f794b6fd42daed950757f5ac5d2ca303e639",
      x"7ead7eb42d46bd736b58f8111fbc1eac0f91927428ad7762d19882462aedf8da",
      x"4851a50a01aaf0ea1cbb9c945cca53b2718556fe687429246ba9a77facfacb8b",
      x"5af275ea6784361d60dc75a193388cde3a94341d26f32bec6983b69a4dae2f02",
      x"f4ea5fa9331581f449a9c4cdd53294ecc16f0dd5a76b75638fb9822d1ba46e18",
      x"1e7863a3418177e1a5a9ed0603da0052a70f87e5f538000e0d922ab1f1561021",
      x"69749ec04081b70e5dc266eac40a63129f857e0df2e151c673d78181e3effdb0",
      x"b05a2216f3f75d2b5e3a9948e986dd02af169c7c8319f5aba7d2730c57a6c42a",
      x"9374f0d5dfc7f2ea68398fd7120352a1f8ec1880e21f7d95cd6abf4f332cbc8f",
      x"f798067862521b33d3fc02c9ada8a59f921460b683bf4f556775a20380578277",
      x"b221a29a9314a702b486f4ab0e84467712c718751f54b9914767521e66893fcd",
      x"5bb9e8c44619ee4ace310e7d9366c7da3c6c379e66aba1eb1077df989d28bbc7",
      x"02f32ce2a965d5d3a2485d4291149c20ad89963bf385d5bbde05eec91de522fe",
      x"73d78621ff81f8f40dfc9d58c6b2477b8d99de5077eb7372cc4a043273128b7f",
      x"397e122c24e7ee52347eedbd4eb9a092c9c9da9414e75150f2e22fee644944d5",
      x"fc1e2a5d8a031d87112efa103e085ddb2c2b82ef283a8bad49a98c0da754e1e9",
      x"7db391a39f125e896a009de0993cbad264a10f3828fa435bd68ad9baee084bb9",
      x"b9c0bbb4e0833e86fa98888d671808c831bb3769a8b1c8fe6ddb0d19db4c178c",
      x"d0d7d5b15f70155070dccdab5574ddac32eed2284588f399c07b5d8ae53ed7f8",
      x"8f4d9cf63227e9bdf3614654665a218f90f011268a0ce93013720dbed8b14f1d",
      x"f32f97e57618f37bb06ec58d91a9b2e5d08629894ac29c56efbed08598a17094",
      x"3a887024e9a4b7dcff9c541d3f843fbdd0b2f4797c32be2f197507abba16b2a6",
      x"c3b0343736d4135fb53553886ae1458d3fd85aa66bdc59149dfa5bea1345b488",
      x"7a5da86422f8d4a15d372a745840f2f638d909e971b27a8696a6e51529eb2523",
      x"f2457cc62deb7acb9c7abb580866c3dde0c47365ecda84599b8a509887fc259b",
      x"7820e0922b70be17270c4d2b083ffa4c8d0e57da0dc039af3a7d540ff8aa69a2",
      x"1192c123b009c30c53a9dda7010bf753307d7dc3824c9ae7b2f8c8949b622bb5",
      x"55a9298805c6d11f09dbc93265a834c1bd082ab38ec9091898d38670179bf691",
      x"2b5635de5af11a5419333a66ce04123024e1ede6298781f7038ad138bdad7331",
      x"b6491aded1c367411b77e215fa87bcfbd47f70e31fb4c8032718810b4dc4d969",
      x"aa4eaf7e6d91ae8a196b9b2f52235e15e9a0eaf966f78b5d2f3b2c1f4cdda34b",
      x"73ede0474e1cbdf031993dc9968e237dc67735a9796cd9df0887e4b1be62333f",
      x"9a3d9abf51a2ef22fad113bc324c5d8c68d433868625e3cf232a01c974f60327",
      x"fdf0e00d410437fb60ea23aed0719dd3cbbab32c0103b45a51fbf267d5c759b8",
      x"e8f0f9065b84913a0da5fc9357e830ac4c7328fe825678a639fb9442fb5766ae",
      x"e930023fe1daa33e0178b1b11daaf6cbe9442249811a61a2c8802fd555f98c5a",
      x"1d1c8a5e9a239044acf85f61124debbf190c5c6a85f5dc7ba7a9b255c53d7af4",
      x"0d53672941a259667661819cf575fdca47b374da46e0d7fd4ae8d3a364233b30",
      x"53612ef915b99a475819bac78b2e15e17d94156fb11e54d446af642835b0d142",
      x"05f766119d68736dc037876adec0d42217b7d57a9fc8cfea1b173cea0e1351b3",
      x"891f9d3ce4388f78be186fb978cffb36c14645483e38fa8c003e3d43ffdbd52f",
      x"bb9700d98d6dd7a1501b99f2fd9e4f77a44d52a2ebb73d55a49d1ce5c342cc53",
      x"59d7430f9907d890a6b0e805f34e54dcf7c84065a6a0c02a51663b3f7abf2ef2",
      x"8e3e1f6f83c508b206ca21c0644fb16c032544af4210489cf9a58e53bb4f1e8f",
      x"b571c3d7aae35cd8b287392398afdee8ce3234aa2dea3785b5c390df7d2ca2f3",
      x"02a3d32a6af929d2798573591c927b0bf7c127f7ba43da82179668aa079f266e",
      x"416cddd788e30712f02f34783bd97ca90625d1f47aa5c177c681135e09baccdd",
      x"0b563c9b145cbb236f8620bff80742c4c95af31b8848cb46679acb1b91df6b0d",
      x"0ef48935e45d6c5625bcef9f856eb75b2414bd1b4a86a4b9b5169fb249a528a3",
      x"85c0e9c19bfa2f798b6aeffd9d84ebde1a702003a47a8358460e66e3ce000b02",
      x"8db02adbaa1a1a0640ae43e27b368b3250152680de465b9824bb0f6a698cd0f4",
      x"aa68811258eff86bdaaef5aa996c32e1bb59378c19b655222a50dadb3723fd3c",
      x"f14b75b894f34184e420cf9ce0a2500caffabc1b4a98046f5517050c4cc2dcfb",
      x"e7aeed11ffc83a73ba2228caad8e3cdbbd0159deff414ecc180bc62e505aa192",
      x"612ff3dcd8082ef959162f1122dd9e38bf30537147372255dab4c34e694b32dc",
      x"9ca7bd869c86b680ea9c9a83979d07ba8dc952367704282a704cc4466b920f88",
      x"6317563cd43e1d50aabc1b48c9d08d1d59bb32c2dbdb2808a107a45acaee1ee3",
      x"10cbbe8f9b6a8e30adb7df4da7301b209633c012b5f6b39471457adc7da798d6",
      x"1e18062aaeee9869634cbdb093ea3f5c6300ef8bc9d29e740c825bb59bea3275",
      x"0a90ae9100d543ee27fc3d77ff2592ae0cd15b96f4a0e953adde812229f9b0cc",
      x"682b5f46ed5783fa279ffaefd8c4978b525d38b6fd0dd92c78fc03cf435bff9e",
      x"f98fbd60b29ad3e3484156622311ba204e74af280ec2980f5d0dd92660cae053",
      x"497ffbb2851a519f5205476cd66197fdd68411e07f0360b70d10556cd8861dc5",
      x"21ff31b077973ed991643c4a1adcef23cb4f82ef91765b800f19de4b70df271c",
      x"1968d76ab25a642c559976eab4ea2c8536dc4ab1bd2d01d19b0368224ab42845",
      x"6f6bf4a6c66b70989578919bde8a2b3402f2a63139806fb9cce8a19f69de11f3",
      x"a83cb1b7e0db0300ac5bce11818b7ef1cd89bbda3ab9bf14d3ce8848a178b734",
      x"ed1a7dc8531ad1478cd0769933ddb0d07d773b47dead0236696f01b3d423fd04",
      x"60d45bc3827bb368e28fdc8e56773d948ec61d5a54a69dd2847cc03b51e0cfa9",
      x"90ed22afd844307273a42a487bb9497600da6476eb6715023722dc270b3e8c89",
      x"30af9ccfae1baf7347c687151e56396718a3d5433e18f62e22e4e0f46b05e8cb",
      x"88589764b906e8711fc33f2fdca975955a16d97fc42273a403a4e9ecc5af034b",
      x"ea3b2360ea309af860fe01a91d94cf60d7b595eef010787acba17046693af597",
      x"1f520052f729e1e63479b23d65c8dbd68ac90f703c3f25dc0e69915e18749925",
      x"b4095731746c79257502f447988786a6441db0a33891363bee73c5eafe0b9b0c",
      x"81ee3a3c51747f27bd57c78b166d5836571435b4ed26e5563bd4af441cec5b1c",
      x"21e6b299ae8ae1fbc0ac7d65652987809759c10ccf22bdf2041b25264d26e5c4",
      x"55544f0b1dbebfc798614bc84480324f77081b1007b704f510f2508613399864",
      x"fe1e600576be6ab4a38bc12c11f33645c569f565cca8165562aa1e685a5034a9",
      x"c948e24859380182a0660c011b136f357ef7b5355b105790bcc03b351676b7e1",
      x"b1f8fdcf882e6737597768cd3c85dd300804a28c232bd6c2033cbef43c3691b7",
      x"6ed5476bf67de705c7658c03b36b9b73ebd70964ae402dbcfbd778adc54ed522",
      x"2e3c1a05ec74e0a6346622b271fa23b2ebb924da07162cfffb8293143edc18c5",
      x"371fd3e089b3e4c9c1bf8a63c210b34324c32a53832e0edb4cc2348882b2c528",
      x"4fb1cf41d41839e19b0c7dd319ef6e3fc31f1fbda9715a76a85365337f10b7f4",
      x"cf14bcbb11aa1461ab2be4ec8f79402268d396b9e3471bc6e3880aafb43de84a",
      x"0ccc9af4226cf85296d0e7bd0a6c2039599bc18a62af614e55cc7e01e322d889",
      x"0265145a29d67c7fcf0af861abf41a15a544f53059b5378db93a5cdfd2e75ec0",
      x"7e280d145f7e0f457eef7188d8cbc4250f6e3043a26e33a43be142152a5a280c",
      x"b80433b672cd5e577c1c2a02f1b5fba503d01eb19ac8710b15faba8acdf15a4b",
      x"c0a93db2547f6e534f6cf781ad1fcadb08b4c1152ae4f9a22e78561200aaa927",
      x"14748261eee7ff017134cc5389ef2977eb08deec1e4cd69b0bdd5785fabc058e",
      x"2188f184443335d6a4a51da7e57d4a6509ac7dfda5e3587568bf1a04bf81a01e",
      x"b0a9a7018afe39ebcb8875b17bc5d6b6b275631a1a5f4aa14b4ec594c2779fbb",
      x"27df7ee4b33454b92a81288c9e8179c6f5115efa03e0c1f6f36809cf5e00a5ea",
      x"f619ff5552bddc2d55d1bad6c1ee55ba01d47e6f81c1d1f46c4c8a360aacb607",
      x"20c220576216d59f8eb24d35c0d6f514bfb9a0ad5971bba5844b73dcb2dad27f",
      x"4f91abf8b1d2caa484e6c3f017c80e31eff8d6c5f0aada36cd4320620cab5eb1",
      x"748b8bafee6816e5c300bec8ce520aa020ee356db7c444ddb6365ed5307e4f1d",
      x"67f5aa3dde1d55d4fee429f8ea65da2ee776ec10a1aa4bb454e019b50e4106c0",
      x"83793c6f8fe863c9d6af6b8df00fb51d22c446fa6b22445cd98453de310bbc80",
      x"0dd3fe2cb900394dfaabd69413571f2d530378b902053f48c44a91343ef8190f",
      x"3848be5eaaa50f757015426da48a5dfc97c45f152f3acda387db7ebe57efcc50",
      x"7cf59e00ac657f48b5ea977460381431d00f3e3f42465fa6acd09f47f9301f3d",
      x"3cac4d3677766c3a73b307ca04e9343f298a8d8da431f2599260f2c83305a0c7",
      x"2a530bc5268afc39cfdb268449ba81978b8085a3c0a7d89f9a7f69d6c4f7fa8c",
      x"6e7b7d387da6f9b85bdeb0fb2a267de333d8dc4c7d45d7ef63292a4407d9db67",
      x"f592e0b756db102603fe4b1158afecb88ffa23ceebc4e04c18b3fe0401ae4809",
      x"b5d6b44e4485ada30c79e7a6942f3ca3fc85e2cb97bedd32496f2d1c5e1d3adb",
      x"edb9ad325dd1294606a4bf236d6c1d1e762866ea870114da595ec331b4da66a0",
      x"3ef09f7f572a348a4fc5916859f24fd12abee5ef05430c985e9f87cb222cf274",
      x"7f5595b2a54c9fcbc06b999d15e443c00566259eda7ae241473730c04ef71134",
      x"70bd2db718c426b22cfec5f457ee101917d246eca7bfe8d607b1f4258d36a242",
      x"3afc6f323afe007f6cdb08591b618d35fadfeb751ecef77417504fc12d4fb065",
      x"60d774100b0b6120d0af542b712321ca79f536b33d3174a8af66d0e951d93f22",
      x"b134bfc37994aa37694256fbdb3e5f6131963e3a39f459835c1a92cff40b9182",
      x"7ea409b8c4f2eb0e927153d2d8eb016aee9f674db7cb2b3091c9de7eb3f4ffc8",
      x"10c53323d95f640a01a3d82698101792797df02048fc40ffd3e75f1c489aec3b",
      x"b2813c320d1317fd795de01786962f75781584b8c46f69980dd60740d6a1d5a3",
      x"2cdf292a2ca16fa501c12120c4c7d11c337e627681980a65ad53f7eb07eba3f1",
      x"28b5fdeaf4eb321b06652b6af6cdab75f5ea7adf452dbe0a65999fa4963eda4a",
      x"e82e9ea869dc5b16f09bd78d32cdd7affbabd8e448c0045546a307c9650de301",
      x"9f238fe626397a49d29ba7e7af74052dde05d1c41dd2169053e2641ffc261134",
      x"3a63a631ca5f6c2a6d682a9d56b7020f9b68a000808030353acb390633b11ca8",
      x"46c2af8646670d4aaea1172c2506bab0539ca844ffa0d694a1d275c4e32db653",
      x"467f350eb7c6071e1b9a4b430d5a45027be9626b0c4d26ff117ccb48101fb522",
      x"608c31ee9bdfdb69196997ee83de9687189310587870d8338aae7ca995762c01",
      x"fc300b3ade38206c2e1d89c35486e77504a7902f6d0ef1a2712a1a393c86c79a",
      x"61cc38aa1bc9769b715be42a2869eea41f633a94dda743ed75a0787e388f1903",
      x"751725c00de65176462c2ada99649149d17ac4ed6944b7f083376e8349a4b02d",
      x"c24f8a973fde4e125ac334ada68fce7ff3c2ae621dcf36c9e89428eaf4f5f5f4",
      x"218ee9bd65ca84c523d6a0543a2fb0bfa7faa151cd07a30c6b27feec289372bf",
      x"f300c8f7d097ab163250e4aea55bc3da6f3a1ad7ea031534210000728c071539",
      x"c7d041ce78fd6f902847590ddcf3439be05dcf030b3227a2375c2e12da698e09",
      x"c18f081782e2dd58db4d70f7bfa06a815e7eb1a73a85f258ad884e15f33fc1ce",
      x"2121cb6a132c89b34f26f6cf0e9d4de05da4185acbdf55e55cf0b7c02ea3ea16",
      x"0068847ad4e991602d4419c55399098671c97adbad79d44c2928b4ea92eff2bc",
      x"f3e1b26912955775176c54f2b88d002d01c71d1d48df40a8c8c6ec34f2b83813",
      x"ea8e94fe55a837e33a6a48bbe875eb0091c01e0658976b2901f525a28101ebaa",
      x"45d61c762b9069022caf77f7722210ad0863f4a7757d2827da066c3ef6dd04b7",
      x"51d8c014a4fecf76a3f61edf613000e55f19686d2e0c60406de91036af40c2a4",
      x"b391d427e0e3b2cd9d47e0995f88757644194288490dad09a2fd3531629de2dc",
      x"beeb8c3ec4eb66e359b090c834ba0405be2ff0e13bb62d989ce513b9f033e007",
      x"d9c12f04c69c0e4a38f64cd155a946a1673e6f0a6f4a30190c8a933040e9ad0f",
      x"e30423d54628baca33a2218432e3254757f3e316ee4e2bd162af696eadaa2493",
      x"1659ee274a9804f1b7eff750bd8c7ebe3315a3f9bcd697195db116d6987fb120",
      x"bc370d915607acc8ae95fa3eb9c00a1896b04e934b96f2cc36b6729bc5586bc5",
      x"402ec45dd90fba346d46fa5c39f4dd819c05db699719e231332bd4607aae2e8f",
      x"7b20ee4a112b9010d2f27f1989852776b5732ad7467d849073f4e6e922b36731"
  );

  constant KMATRIX : T_KMATRIX := (
    (
      x"0d2f5f5f3cfd4463eb86738295cd0f84b4da42a6db04bed6913a373429b9ecee",
      x"c720f317af787853b1d1f0ea110aef330acae297d7c5855f40ccd73cbdb80e3d",
      x"6f789b4e07eb3dff4fd4a902de924ced9aa618554deaf8035e9ab97e660ce1ce",
      x"ebb36404920a76fefbd944f2a63aa33ae2558c807dcc29ca5ce706247c23f070",
      x"cec02aa03a4390fc2bf7c0e5fc2be3d5e73a819bd064a170a1d102206b6e0c4c",
      x"c4fe705a6418e9dfe445736e903c02a6a364d881d9914cf4cd8393852a65f04a",
      x"923481d4ea338f64693065ee03f652511578ea9f0b17e1ebebc5d552b861e2d4",
      x"253531ab5710882a2867589d5fa3ddf9db951ce524cbd3a9bbe590c4663191b4",
      x"b806ae845f30a73d587665a3cb4460955d01489e4face459ccc291f37520b809",
      x"e3666b84ee7f1caae7d57016465dc8521747782b32bc5806f9d8541b3ef3d89f",
      x"ed78860c94c8f156805697154988a021a16a3a86846df7971af85b2bea7e6460",
      x"f5f0aaaf3a9bd6ca7be4d1bcd0e4a64a0e5e30751d5c7f4804b540ab07dedffc",
      x"00c3d99b4378e6c39292feebcf58e772d31f6526642e5a2be079a3797ea4a25a",
      x"10990154edf80eba34a416a0f5d6503cbd85ca2168c2d9fa7baea7682e6d0d33",
      x"aaa67a26a2c81501abbde83f1b5d941b245af57e96637bbe2a6c2fa097f86eab",
      x"5f27de53b4c30557bc9f0c833f1466938445ac4dfa5cb52e28b26de77b80e6bf",
      x"2e6c855c52924d0bf6909adf5f55bf807ba45c6610136d6ca226b747742af649",
      x"54d3ffd883ef6fd17bb8b257be7536161d8a8d15b32eb6397994d41aabbe8c48",
      x"2c38134fbb1a16cdf8f9b0c09454f9f66cbc9a32fd1c2d1f8e44850f234ea1f2",
      x"50794ece786fb5083851b2cca385961fc20fd429b0c2883bc837e0215ffe6e4f",
      x"889fd409e2fe4cad0d73184a3903f0d2de2e02dc81d559fc8cd9e3b4b4ff72f0",
      x"3a2337477c9a4d64d017d3d56953c467ab53691a3840933730f0130204f26550",
      x"23082485f9fa2a45100b9b330e457ce939f40566657fc4af937a8176f60f9471",
      x"b0bbaeecfe831f1dc005ad9d9ba52cae378a43a61ebed5393e0215175d2fcd48",
      x"b521fe7f11405a656044ab316467b2fa04c660d72419013def84de7e58aaadd7",
      x"803bc6cf273ce8461bb08cb3e528c6618451b73547b026792c93bcbe8d6ef5b4",
      x"4294a49a8b966e1c25eca3413ffd92444833d4a7d7ae74639ab4ad21305cbd4a",
      x"7fe62a9398c7ea5f8219af7136610bf85ae320842fbb64fd47f0266638508efd",
      x"71f3698c23f15c0ef61410985c5c74ea20f32be34ce15c24e0e7f85a56c39534",
      x"6d26345d913c7324b1f27788cfc227ed1547d0bfd711227fc84ca85039ac2ede"
    ),
    (
      x"c27718434c4f879128652de0109ab8ae8aaa103c225ed7fa6be42a1fa20e8e23",
      x"f3a56fb1e72c6edd78fba9ba41ea10cf0491e8c42193fdf39c86b023d6430c06",
      x"ac7d41a4a103c73b104bdd2cef1625b5ee49259a5b866d4327e8366050f27536",
      x"829f29d168bf2997fede572901fd2d2a9d08a9fa12d5a564884fbd23a50902c0",
      x"9736c22e446b92406b3fe90d26b1ee75e79cd81203581001a9e1cf9f5788ed94",
      x"f05ac30ca027a3c7fe3809073c49dc1522b1c189878e4cfdd2be5e04e7a33527",
      x"ddd81b81e2f4397131d6e3bd74b36cdff6b1ce599d4b32ab64d2fe2d38cfdcf9",
      x"62d710c3fff1b5f2693ae50ddc0e96c7f47c130ce4f66b0528093a4d286b68cc",
      x"9903e23b34286c8c9353b1df9071caaae667efb106e3ae40606f37888a7e6360",
      x"09251cb34f6e037fd0e4f951151f81ddf7d9c25f10759badc4c4f9e7d5319647",
      x"e9ed29166558e8a149286be45cd55abc2272fc6ba0f904f50f7b800e39f05e5c",
      x"9125bb2b95a67ec27817cb6969f2cf0c49e51dd9db228944dc20fe201cfb851b",
      x"9fc7ede956fbf4d76a945e3133808f1e40ee3080384e94885c2442946f051793",
      x"a7c595da2a79901ee3d0a4db28570c6d8cce8839627b09c447a1373fae95f0e0",
      x"c783baf180a8ee0f18d5cb476ccd8176bb8c22d9a7ea333d7cdf72b4c38f4377",
      x"f2a5aa5f68e47ec159d6ae1f610f6fec8d5d16952688669c781ecf4df6bfe29e",
      x"3d020713f5070ccfdac7ce60eafe676697deb7d819631e9847656b91405076f4",
      x"1b11f76e64da67a6622ca14675a0a9e67c83f2492020bc9321c3812f1a5195a5",
      x"b7808b4cd7bbb60d51255b74095b72e2bfa1c63cff986f5ce3ecbfcee80d56fc",
      x"09385cff21589396e40ff0c4895cdc8ec445d4f56e9e4b5a2becebf103720ae8",
      x"0e17732fe0372ed597b15c221e869c0c19c4203e910962f5ecc7017cadb38faf",
      x"8bc9dcbc3dae3050514cf4fe7f1389213770d05536740c5ac29f8ca9647ae2d9",
      x"a6c0ab687a05e831b74313c772c50ef9686206f9b10ed0094795c6de892ba777",
      x"c588c44d67d37eab6bc55d0365ac227b7c7088afe4df42bf25379621369729b8",
      x"7e707ef947d8de5ba1731f35606c71385a17ce5ac6498661e1a7941f46b9bc56",
      x"4bef4830d2543339d02092d45418b70e3f1ea27b56d417635be0bc3bd902685d",
      x"60581dd10cca3f1143caf59aeb874cf532e67c8f5ccb28ebc46e791f7284c65e",
      x"ceda940850243d5233ad80a2d65310eddef050321441fddbdfd8da630a8e5fd0",
      x"8e26636387b47de2e91800b10bc3be283f7e4420186bb8eaf8a930580c9234a7",
      x"b0f6a919db22b17e7030f11405e803bf036ca7fed71c036b3e84ff8e030c0388"
    ),
    (
      x"d5da3e32d9633d64e2c875408b990bf07ba613cb8186fd0fa761138f045d1315",
      x"a31226ab2537996fcc8595d41c914e48358c864948edc2653956d6f7e5edc71b",
      x"8fd7af94d00426700adbede960436dd6849d1e362d27c310d06cc5e9d442a625",
      x"7b6c8fe65cfd07f142293ee0e8a0b399691ff0e6287249fdd5672414cc93802f",
      x"9d22cd0b150149ba32cde5fafce4828a50f28b50ce4ed876f4935eaf2fbcbb60",
      x"9686deeb1f537ee21dbd7cd07a2fb7f6d6cb8f20a6a74ff65a149d25d232c754",
      x"6fc89641bcfbdbdf549929bcfed05c9a6907077712ec7745fde530d26d5b7bfe",
      x"8067e0d8597c92744fcab3648481f73015b16911571bfa44e0e79413a13fb421",
      x"0b5f00a205a3fc3249337eb9f87dab09e5fb671daa8792cd663c64d378876fa9",
      x"3dbc7feac0b88154c820775616d55d34c79ad2ada9cf386d50c7446e36917ba4",
      x"f86b1246a362d0b55e042027ae9a4e913ab7f171f44fa9e6cc9792ad8aaeba81",
      x"79a6e420c68ba8b94cdfe7762734878c08f676a3f66b1916fc4939899a5174ad",
      x"02e03da999ef37b9a0617ddbc8400fe1acc09952ccd2ae251730fbf0b29bba18",
      x"4257e4b71a4e74e876669e1bb5ef740c16a717de9aa22f32fa1d7a36f63982c7",
      x"f0399a6c78c8512e200ad550080530404e1ba58fc7c2e848fc21306ebf5d8eaa",
      x"1310a2d81966a9285ff180e6c4f68b3c3c2c292d59cb72e7fea3f998621147e7",
      x"b59c51703527f495216ebd0294976257d1f93c6ade0ea60941bc00e34faf1b06",
      x"e53a17232ee6f07ac2e81f91145f272face5f126697a5ae93ec1c49a444e8539",
      x"994887090e8e6f66559b6118bf954f4da2076380a97619b091601ced8f57e39d",
      x"5ac81ef574b41be010f6f8ee1c0b24ff1a86055db0115574d5833b97c5b00c9a",
      x"2e3a19d310d51e9c246fbb94281a223684455dd6810881d5c5fe8b7ba20fa8ba",
      x"78db86a0cdd66121885e125f43d91b38b935de4c277c768201a44510a93d607c",
      x"e16923c83811aeb8cb54e3c581958cf77b8fa118df03aabd916a2605aef982b2",
      x"0881b1d80f26d84019a198ec1dd8f89381d3cd9d09f34e38f5298f893ce3c110",
      x"354b232d7963557c088094af696232f67eb3c4ce2dd6df1b55dc778cad48baaa",
      x"d89404b80963214fc45577dfd155fff7667596490302222d0558e7c0fa1ab273",
      x"1b8b62113b498767f001fd820597ad199f59e0d5cce39912b3ac60b54a825160",
      x"931acf8a5d1f047212b8f059d0ce7426bfc7f33846e080a9dd189673b1d828bd",
      x"39ae142894b6fa05b6c6172cc6d537310630412ae46ded69fd562cc06832bde7",
      x"ecebf6dd50a68926f6c7419da5b8c85ac102ff99e52d5889f92220ebbe8bd4f5"
    ),
    (
      x"9fad3d579487790f73b773b84c7369bf9955aabb6e186256bfbfaab88baa9e8f",
      x"84a2e73b29dd0071ea801b87160cc40834af443987c939122c438176c4c29c97",
      x"9eb9bf9b9e037e98b48d0a8b31de63a508d2d1ebce806f2b364204bb27058467",
      x"1d39c42959360a120c67c09dcfe7058770fac581e71752c57f865190ab45938c",
      x"368001737035b3f96cf37897b8c1b1cb5aa0dfd0b5980bd15fbde70335e2fa1f",
      x"fda77ccbc69e4f1d8b1e75a9c3b077fb30cec6a04a2ff149028f9abec2570705",
      x"0fdf332c736572a68ae00e3a4bdac22f5f79450592daef91aaa03ee040ee1557",
      x"0c0631464b75e1d506e3acb03ce095793f5490a257b1f64b3a41f855e870aa07",
      x"02041364a007375b225c98a5c8e89c4eb9084ac10e03cdb42a51967e8a6f9d28",
      x"88f938c0001a3d4e40099b5aa77f2d97ce36228ff1fee981908cc94e75f6c8fb",
      x"76ae3fdbcc6d9787fe90ef1a83e6b40b3435832ce51edca637eac7344fc84234",
      x"51c672766b88f73042f1c3afc76c405c3f28c973894bf08ff72ba9d2fc9db451",
      x"c94d3bef04a0f6f603a6f2eb9aa80191af3763330791784273efb1f85e1f893f",
      x"ff4b1d7eeb761c61d4e141811d53faac07c1b408e1bf902e1564ae6411084410",
      x"aea019d2c9497bb9ea2fb9fd555b7cd9870698f5d6ca013ff6cfe9a45c12b598",
      x"143841fbce333ab91c2fc74a90f02bbf51fdff785f3413c8b0d0c2b40815c83d",
      x"53bbafde46793476e537dd75b2a5e791db4f7caa9beda7f07bdc8a6e31546067",
      x"97d92752edc17a0a84ce0b07940d1fea75d3ba150dae7f3056edec037f4d65a0",
      x"949c64264106c5b9f7c7c49e8b627bfc0567eb159600aa0f6b803a962a7d1135",
      x"41d843b25726b17124752e540fd9a925d7d9184d333b5c950094dad72e4adae9",
      x"6299763bb1460e45cff7fd69bd65eb4ae31b1e28c9cded214fe91b8d4ca1dac8",
      x"d7bd89f15495417e342ed9ead343e6203a3571e5d17ef88f0b89ad0b4d945d48",
      x"db07ebc3fe9cdf3585d2696d7c99f6f8c209cb77358bac468c4c0af0440fc0ab",
      x"de549b41c7ada96edf6a0ce8948a95e45a56b726ec7e7ad2c6957e0a14e744f2",
      x"4cc8de3d4a3ce874826131a247ea4ba1668a076e4333a2379e12ba349dffcd58",
      x"647c97d2b551f0019a7ef48e623c8c060d77778113da22ffc06a2ca1cbf8bd99",
      x"98cd6f57ec87d8176f90cfea203a6655710b5efcb2c0ce79688d6b38b7ff3d4c",
      x"4ea4f87e0aaabbc10f03828ee75d0c7278d9bf8c0c03b627a99a78862684f051",
      x"8ff64104262820e4dee0a086d974b683274ec6f2b598a226a4a41c0c8a4069f0",
      x"5a55f2592e882b3c6cea17506816ad2d62088a85d9a61c70ae392b5f8c0c1f98"
    ),
    (
      x"2665391e672ce88919894686f9629ef150723865fdc3a7978d1c6a1f5c1fc140",
      x"ded66520ad5aaf0160915abf3049ed19459dea90de3f24d01cd544a5be1c3f3f",
      x"0ac0a90c65df3386aa72fb1b811e58a8a0ad1cec679a4b66103d2b607a03c275",
      x"0e643725be8ec4872eab429ae5229c46d8fc64c2e38a4a176521dc1b54e0c03b",
      x"baf8d9ec280b85c0a3c3104171b1c549c53a7457c190388e4142566cbd9428a4",
      x"447b3343ebb5dd69e8c97f8712a7a9351aea5422df7ea2d46bf5d0e2f3a7552f",
      x"43c290725002227d4bc4177fa934868fc80189b39b051376f0b7a925bfcbbe14",
      x"5dc1ccf2b2c632ba1c06baf50dfeb6533dbffa1da6fcbcb1a33502f07f9c8a24",
      x"addb6913ad94367032cde9c813bf9460fe6434c7d7b9732e13b25e065314e0b4",
      x"9a30ceff9e022f8329185d3d419d8a1b501d3fa73b981a42a397dfdf576f8b36",
      x"9edf7913e9fab296f4bb867c6ead4c98821734f8a68c05d49043f4508f891a05",
      x"b54d1f0142f3d71020a8b4bbf4d66730df9952fdae2fc4e28b3d01baa79ac427",
      x"382e5f56a158097f193807c656170d9b89efad2b6bbe71e6b1796fded97ca20e",
      x"18e4e473fe95e8ac8ea1a380f3b09234213c32f4ea78bea2466576eb752ca241",
      x"92937def14b3ba56a261b70114386d7f564143315e0e89a664c9ecd0da98d291",
      x"bf51d6ad3100c2b52b255dec347e2a2b3aa7380fd47d9b114ec08109de74946f",
      x"ea3f68697dfcfb49f1998dd2788d58fb0436ea075b1b43c783474fcb8bbee7a4",
      x"b1976baeb39b3d31cd2c674e366f47831f251de0c1850743058e8f32d97fcd27",
      x"5db4b214ba7a8796cc305e1d6dff82fe0c13ec65401610676236dabd6fe6c3b6",
      x"be571dacd82227fc65381ad73488b66d04af921d72c4163cd1f08dca8f5fb565",
      x"b49a7c49d521534ded3e48836611b554f00549440c74ec6833dfd366850d9f87",
      x"e5109abf19688923073b4664ea795cf06f93c7d2f8122ecd0c88a7e2ea28883d",
      x"ce08ad9723121c54f38b05164e22c69d0ce1f594b49943a9624bf7cb8132a3d7",
      x"0bbb65b3441da2146a2cd203e45d7d8bb7b9ebafae6bb5346a226a5cb1d492dc",
      x"4e9898fe4aacce3bea56d48b9041e15bd89f483ac1b0052cc2eda5e1390fa22a",
      x"48321d29cd8a3b4750f778bcfacfab3695d40e690730e41834ee7dab05e9d494",
      x"b2a17a7ae7ffd9c84ce0ec6014ec41555f657947fa1bd25444cbefd6cca598df",
      x"791480bfa983aa7e58a88ebfb8e88219217d918b6d3431748f63c1564572e158",
      x"559e4653c9b6ddd4d0944b05029a66171b07ca9347a15c49c7d032dd7b0da7d2",
      x"6199c5288478d4fbcc22f5ca74d5cae2cd73f73ec19e533a0f4464b670aa4447"
    ),
    (
      x"273be703a31223440066fb7a9f0f0aab9c2805311cbd974a953d16fb316d83e4",
      x"e7e440dd1773dce42b3cfd2f7057704145b334070fba7558ad7545acf09c6eab",
      x"08dce157cb5a2d6cc48e6a49a8c95d8892cefb9257ff3dab734fa877cb228c3f",
      x"64a3132754a6032c652dcca2a0116164b528dea918bf06dfbe518a7334878d5f",
      x"71bd54dac5447fdbbe5d5ae0a68836a67f17eaa9f6b7f15143131c1ad10c8d59",
      x"e254c7acd7e9671f9257f66c3e1fc2fd098eb85e014729a2039899ab8d128092",
      x"f140edfa8959ceb03ef7f7f334e981ae9510e0fa74de1df2432147ed5565f9c3",
      x"fb094feae09d21af5a1d34bff4a6f2c099332c98bd5ca525136114e90751aa2e",
      x"a7304899329cf668c0ab4bd9b56b24f0269b8f13a35281ee42c14bff34731799",
      x"7bb4fb063261ffe2d340ba9370d6029973e7f50d98026dc4a26742c4210f8501",
      x"bd26ff6b54e5d1ed52d8300e960a9ffa17478c548a54ff8bbff03f2dde57b687",
      x"0d6c152effd09659b9fd30123ccc9a92ba02852268f88a29b4d2be5c9743a51e",
      x"703ccf22c11c24af2b4bee6cc8c88467cee568f9aa5b5c2935392fee6917edc7",
      x"87dce489849b434f47e2e0f904831527aed123d750a5770900aaecf676fdafb2",
      x"38d5e470da8ac9c4615e61dea29803fb83e0e4951d786770ddd54949b55735d3",
      x"56def5aa292a1360802a8499fe1673705362d6495058f329a28b079c9900f24b",
      x"b8f393dfb28099d5b5b958f67e0847d39b7192d4238139cddfcbc4b56fd65cfa",
      x"df52c4256d42a29015ea1f697855d0231e98d9b5b919740f0679c2a928312cd6",
      x"5f75ff71eae05800b1d30785c15fa13af527a71ad3a0dcd94691e6d0b5aac6b9",
      x"335d3409f0161d6ed1f97501f6d24c269760cd61514262779acb87095b4ea62f",
      x"5e1f10b3dbe94eaca137a87364b5a3e382a80388937acecf5ded99c4f25ca756",
      x"6a87061431f84c873dc72548ce4fbb6c5c805609ef60e23fd3d2cd5ad6ed9fa9",
      x"0836cbc2a06f5283350e896293a795511dfdaf19b7480ff7ed2c4705726a1da4",
      x"c4b1b6460c8784b0654104dca1694cd7ea65daf941d37dc8bc539a21b7cdaa82",
      x"74ee22057204295ccebe00eed1e2de0f836dabd0216437e7b644c56658adb17d",
      x"dbd7c0a0f44bd5adfe309bd67e9be41d7c4de57f27d0e95752d36e3f2529aee5",
      x"aeffafb01862eb350fa1bfa8347cca8324c4d6137a1f3e1859c9b5df4698f04e",
      x"bad19ab1b180b63ec4d4b01de442fa979a383441b5857cfcf94fb19c49d57b64",
      x"fcbdcba52e441e200205dc6d61e96dd9b5771ae1ea5273b0d4f604bf10d19721",
      x"144200a7c5dfe265d5a8a87a9369500bb956d4984d1c3db69e5950d795be1187"
    ),
    (
      x"79f3258dfa3408f9b4c5d64625c722f18c1e553c870f438a848b12c8f391b07a",
      x"d967a9dcc177b9ae51eec39e4757679ce588f2300c92e459c83a679744d672dc",
      x"9b37537b2b28ff89cf3ab52a1323a21bffa85d9e7d283ffdeba7f1327aa66190",
      x"924a6799020d9b76158fff3cb81bc9e6e0a94712166f77d09856bd89a4b6f50a",
      x"4b87dc399809df1acbe4354f384149bd8cd5a8b9f0c0191a2eb5471f833f1bc8",
      x"35d9635db7d368bae649bff508b509fcd937a2241381b33ef0fddc5cc742d9b9",
      x"76860ee6081cb8efd1da272a44e6b4554e7b65b09dc1fa2e21aa7e766b727840",
      x"4b4d925048362ed0dcd4016a631d0a109b252e78c6c58f13e7438869fb0007d5",
      x"8f71a0aba5be57676be5fb872a6bdd59b766933d185b67b5933216b0a39d72d6",
      x"e26301b9a923933ce4d30f05b0fb3664a0ab1b14a6f3dfebf6aa77de782fac80",
      x"38ad40b6271058a4e81cebda463c7277eb9f7183c79ff33424829f6d8fca3267",
      x"f6b1cbd6f7168a452a9ae0a81adb675d88d792d10eb54bc0befccb053274b273",
      x"88b5cf45df62ae73394d2c90c1f57bb9f11f989fb435c1cb75f8240c792dbfb9",
      x"993a2a3bb554a3be57c5b0081bebe95dbbfc46c77644973c1c4b6b9e968c0eb6",
      x"53a08a4bd3bdf0289edd8dd435f17a7c2be0bb6161d3f0871348ea7b7f26a9ee",
      x"eaa3abdcb78ba5b754f5a8457050f149d40f6bf551c478c9e8d43fd469b39ef3",
      x"83ba3f4d7a14afab20d7461499bf10c1c6832777727183a759d4ea43b6d57c11",
      x"7eb3c94dcaa129e49fe147cfaafca5e3c51a0946460eecba8ab90a69fbdce42d",
      x"ef262ab61cdc32b466b566a50cc2b671d55d056ea2ed2a4715ca7b8e6407ada3",
      x"9a8dd7ea7388f23add65e0626f04477e7b8a9bd4c5389a68149d7c16e1348c6b",
      x"7f706d7492718ed8c1f081e63702e99744d5541f4889ab19f51fbb66272bd696",
      x"793f990bf3bbaaa95c09f553e7c7bd8e3c18dce35337a1062bcb815483bf9e44",
      x"6cc9e241da948e0da757e970fe58f7e82729e586c1514f70b670b2ce6b402e64",
      x"8650c99b4651765658c6668450e5e4ca56a6e58a6b10e58063d8852d30eb0c71",
      x"2168ca131b6f2c088539292af9d1945da66d9a3daf38ec5e79a2bfc240dac20b",
      x"462e3a6475dd3bd460c36bb38b7e4761eac989df1f3fc85f2768fb46cc2218c8",
      x"054943e8ac094ee8df527bd8bc87cd16a5159332f66771ded50452b8ca9838c0",
      x"a20e2b837dc78b12b53b4332c07d11f67a93d9bffb3cdc44b4c3f84c2a9c00cc",
      x"680a8cdf941b6e9935737014e5893c9e8ead0e9f4bed3ce8138ad22a5309e21c",
      x"9e0d7d23e5d47bbdeb7962741bd66d1131468738aa4558b6d03e7cef8913f8a2"
    ),
    (
      x"b3b3873a8ea8d6591f9eb557d131674e5f9ebd2312f8df59605c1381b0232c5f",
      x"18e6a2ad9cbcfa0abc30462a2a26dba5f6c8ddf34f81c67fb7d41867b0fbc3d0",
      x"3904b9887fcd6456550c2e5e966d3f66d2ae1bc4cbb85444a5630e7939e28d08",
      x"333b52e5ebadf382484823fa65a34c7923e7a2a4faabafc7e471cc53ee86deda",
      x"6733362e3d6013dcf14b3f401cb666317a06f99af7f49a8fdfb99fd0a1b66a7d",
      x"1184c3cda0626b9b19ee71eb268db6ac08bdc8704341f971c92431f176551aaf",
      x"a76bdb0d054980495633a074a4724eadf56cd090a78a09a1973d3b3a11b2cf47",
      x"b0b7c8fac6562a59a1fb49c6584d6eea5d1141a7f6aa96df10d360f82df37d46",
      x"4189c725a97d67df715b111d9ac39ce4d4a234d40c372122bb78a350f1add4ee",
      x"580d6e36abf2bf97be6d4fd8b9e6d3355e63911814f8448a928e14ded2759ab2",
      x"b7b210c6f8b127f437b0b12fc6bf4ac88ec6fc283d7017df82fe4431b5f811d3",
      x"645a2ef598ceb79ae69a5b096cb8e3412408822f3c57e0f1970e359cd520707d",
      x"477360c48caefd568c554d574539b3b866b0c20fbcf4463ebf4b9ffc74675698",
      x"7ba3d74b0e447dd24730512a42de846031fac4b7a412fe076104a02bfc66233c",
      x"9e99b0f255454d6bf7b47cb208e6788abae990ae4194df13c77330a2a720b19c",
      x"4d08704b8b026716773694e0be42a225c3ec650183ae351c8bf3ddbd8ec02120",
      x"5498f7534383ebed25eaf6c31a7d4e88e6aa32f7e938d759bb53e2084def2316",
      x"132cd43545d7c5d72f9f0456e94b28019fc32b2894329b7a75923df74d8462e0",
      x"8b00c77aa01fffd94ac5f132784d1504d6869dab4268896f826b434909098519",
      x"b13adc51d9d2b58f876b43445b1fc72b83be18d8f4702828ce64817f3c249862",
      x"dfe23ab641e777b8d2848c14a02c49155ef2fce4cd164543135650ff541a0f88",
      x"eca5a43c205b0871c3a4c9c7dab14314f9d5c35eb8d4aa2833a974a7e6313c0d",
      x"9c9fac7451721b66e38c54fe28c6e082ad06130765b610718cd0e5d8db456c17",
      x"13400b4077fb61357c0c5d4e186f677cadd0decf73b13c919118bcb056f345cc",
      x"2f8dbe46df41d63b86214cc352d24c8e44648edb5bae8a56079987609f9e005d",
      x"c474a183494b34faa69dbf39017b12b3e81bffd562670b538dd4b871b2732c98",
      x"5a98e8b4518588d606ea3f47390568de216370e427885e10ee974daa2ec82021",
      x"d5aefba35a054132fa506ee731a24dca0e6661e55b86b10e1363576683f36eaa",
      x"8526537e3933d66f6ab25033580dac9940f3069be090615af461590aeb90086b",
      x"6b71fd6dd8b2ea9c6d447d37193cbbb578f7587cea13ed36e4a12f89ac22a1d8"
    ),
    (
      x"0f280389a381ca0753eec0ce0b6c3ab4078f12ffbdc57230c577acdbef9441b3",
      x"0bc29bb0fdaf4a012c06280e5306ed69962c6ab0a57592d12944b8466b9a4c83",
      x"5923062e45173aff001567b10cb1a1680e80c2ddeac7ffedc1648819e3636bda",
      x"ec19b80e0a4e09e90ef1b8b56d8fe1634844a1bb7ad27c6c6e71bcdb5c84f0a7",
      x"723442686ba2335a528c29083328d374ac6f8fb84933879bcb1f7db63eae9d75",
      x"f6bbe331625c85e881b444acdace6efdaa5b923e2ad6b5391f533ad0395deb45",
      x"98d837a11ff99edefa030dba4d7baeb7929dd9e24ae6ff7f90b4440882f6deba",
      x"b2b2af255bc82f75305c729c20f85238c0a7db890d0f7f634d6c489a36c14b5a",
      x"d44e8fba934dc433d7be6849eeda29d437be5cab62c4cf0ab1a7e4aa7d3e782e",
      x"46515b895f97360421347f526a68eccb4c926c0067b2fb5a1ee5b33d944b798e",
      x"b35a068fdc6da09e3cf8e870b606fddd7d786e102f354887f9818a1c4d45d736",
      x"1434b9f8f6dde03163014a80a61515f877402fc53c0dc54b4a1ba267092550bd",
      x"cdaff56693d85c81457d0a5f091b1f223c06306c0974af130db7e5dbc21f5a6c",
      x"a3c175d0cd5a2fc2cf40cb63c1192a9c9c3c4c8e8b2adede39f70f89c6b765ca",
      x"7cecb817382f92a2f15f1fc1762e95e23c088c082782927971f76f0f71baf8b9",
      x"0d74d4609d33980a3846620aad918ba17b33d5626753ed48014b576ad84fbfb2",
      x"76c2856dda2dd6e04a56afa0b9e97a9f351c86fe04e44d131a6293686217d7d0",
      x"daf5bd6eee8367071ce4272d765fb864b8d7ed6ae4011fd64d13e1779337ffc5",
      x"56e9f2359b185a447c7c82288997ede1133fe612f953e9b7b5e3cadb020a2cbd",
      x"45e3896b36c173f74a6200f7d36f0c76b83bb1bf9d9b91ea6a91180666455a07",
      x"70e13219ea3f772745e80a7d660e667c293914e1d587b57f1098c8c6eabb56ef",
      x"48957c5373b98503191e3cdf0dd7a0d58a54a38afbc7a3160937b0c0d302ce03",
      x"fdc2200e33657701a649e4d5230084fee4ebcb8cc029d5a68cf43f81329ad4ff",
      x"40d19064b8ddad9ac391a0b3d4c87b897f96b38eb38edacedfc327baa1f9f92a",
      x"05a2dccba738d797d7b4a98cc323b43b5c11dbc332f1942af0ff4495385b1fd0",
      x"4d9db905cb714a914aa37197481f8f4386c7474cf366bc8290ae04f498ebdcf2",
      x"dac0d1b56d498d472c37beff747e001a83a2e96928018adb33fc8bf7853e8d4c",
      x"f8c1c28cfd235edc7e7609e23e21e9fbd79841bafb4f1c6f1a78d62eb99e7a7d",
      x"8786eda5b91d6701e83d4428d0848d7263e026576c466ecaed02a2ac04e651cd",
      x"5797864636aef76b6c2338761238c5e443a29e454fa92e4dcdba4645eeb5ebbb"
    ),
    (
      x"98036eef969c7d99c2fc73b9469d5b8f1152aad1056c5349657c16b105f2eafa",
      x"1b383bbb1de30c91c30ba0d39b0195ed9403b81223389a9d5a2193e84b61b2f1",
      x"d20c9be3272aa65a35c6c4105a97f30c8e181920724e5cb19ec948030c2c2bf0",
      x"f86b359d457837c9eb7611d223dc9b628ee15d3fdb46ad4ea1896f5cd1a826e9",
      x"8bc57ae4bce0c776ea71e9f4e0a68986bf61e190ef296f25a5f95535e7aaeab4",
      x"20ca27b6befa94c81299f7d36d884105901db457c7407f074babc1340970a7de",
      x"f66a5d7d759fc8eaf7708a4fac93132739992cfd208f1bb95af527d4c74cb87a",
      x"ed3baf6ef1998cc69ff780a622ee507804895f51cd6222aa55eee62d61a72892",
      x"97b1f0cf6f9b20fe0ba5aa13589ea45f05114ab164de1b769c162c05f40b6698",
      x"9fcf3888fbcedeaa7f24112b7a357bae238805a2eb5fa5490d03b884e0b9e490",
      x"4cc55af56a7d298b314416be3ea63b133456043c427071441dd60b61bee929d0",
      x"eda29121ebd0b8844a31b6bf7146297876d35dd5f5a14c0cf3f059df7cabeff6",
      x"c1710650f57020c73d6236872fe722405e85d8a1e8c7be66fd85f2bcb54d408a",
      x"2397019d41298bac564a953cc622994a2e4831298b41de0669f5a8d0396b4ea3",
      x"ca2a2f0af65639bc15778bbb7c257fc814b8727136735be7e18b81cd5dc461e7",
      x"fa745a1e1d8e1f7ae3487921df9576ba58b7f82dd3a6d0d6a3f6cf3b16ec68f2",
      x"7b54e196ec08c58c6575d123ec28ef685c0ef4462eee979800e1aae154c6f6a1",
      x"3344a8c2b29eadd28711b887a024bb2d9922a284c1eeaf86824bc8749e401001",
      x"f0d0f9a35d1bb3ae63f9b9f1e19e18f9b82f22adaf8d1ec7697eb047883838fe",
      x"3fb8f6c2e065a8847b3f77a42b7428c7b20dfed71d95733bfd4c71219280b720",
      x"f11f719c6afc437d6287cdec1037eb5e409e777aaf51b5e8ebd1d7e7542de406",
      x"d567b9b5db955af1acb5913910ab25ae78c259b86d11174835a854230eee0cb5",
      x"139bc7cff4fa5773c4db495dac1de8e43854897cab4e78bbe14298cf48638c43",
      x"de3529322498fb96d73cfcfb0195698764222311d0f1ee5ce5faffd4b13c1c1b",
      x"b09b3753db009924c73366a0fef9322099b87ecc93c6b25dd4f01129f25809c9",
      x"6622e0ba3274a9105d462f9034046492737b833d2992f64aa5381eb8b443d4d2",
      x"7bcbeed79880f44b38edf68be621b22d8e17713ed5fafc906ab9b33828f9fc79",
      x"7f7815ec89273cc8e0b99e01d082ae45f34c170ac28e85a3903106b7c021e154",
      x"9039908d890aad5b89f030138ac5c92e584835af277e3cb4ebf4f63b257e3d6f",
      x"90d0041f934966fd760eaa274af84a7cfab03176301748e786e245454460e4e9"
    ),
    (
      x"b156a80739a5dbec08818739b122fda03c4c34088ef0848544b8a591b44b4080",
      x"044a045de1a3a504acd40f09659ba8ce57f2bbc940d69521e64d61fe4ef73efa",
      x"3819b5e4cf1fa7a83d84141c506cdfbee6f20c8a8e619d3e3f74c6f4da634ec1",
      x"f622eefbb08232e8f9f0f0d6f502520ac1fb6280d1d94b335703833c0b71230e",
      x"c5c75ea7c748b9aa964560523b4eda5cdd095e00a4c95b99884c813e9701f741",
      x"b7e690739d76641b55b724c5819f94cf7de21c1ce9c4f09a6d50e803509085c5",
      x"fc0ac3cac393114d68e830c8bf9284864eb8035da518c5c4403cc8683f0236e5",
      x"cb7cf306c4c2b7876df8c2f64c6ce48f3fe58b56b6f45350a9c366fe7bf5edee",
      x"cc76887d601c3d40a44f37305912d2ab48c4af97d691bb9476cf7a336fc25a9c",
      x"2afb4a809225da24e8bdbbddb73804af443b1cf335c9c8f1560a08e20c62a881",
      x"cbab2ede12a424b3fc6e92f287579cf904570fa92464a8f73c22f766b382b4fb",
      x"9350571161cd8734561616b00dea264c9f6a3e9053ffcda4e5337ecc27055d4d",
      x"7ff04c5be327bbf9e9e67d83d10f0a1052ef1e0e8e9e9da951ecdb6b4492af3d",
      x"13d6f4922e138142f5dd38644c6d46abac1a81d333a1b9c782c30e0e2ae75e3c",
      x"304b8f2c1b1c4e56ac74e5832523345b402d3a2f8715ee79104e25a6e1fffad6",
      x"d3dc89854f4a15de2cf525d720feb40455222515d59e3e1ecd5d67c94978adb7",
      x"426dc7e3c70fce5068d48a4227e64a65eead3065d1e99e0b5d572fe48bbf83c0",
      x"368ea85ddf53933c6364186c4d45dd8aada4e8989d522098e6a34c5517edd8a0",
      x"de7ddb7a6b2a40a7e0b47a5a4a8726216d32cedb4e7ed541fcd49e101cfaf29f",
      x"70d46d42b50611f394f3f1c7790cc7e08a832e6fe750ab88ccbf24325b0b5aa2",
      x"7ca78f9781ccbb0bfe99cc4ae23c52329338d82e131d344667e8e5af314e6423",
      x"5ffc34ac72a5f246794ddca4cae166ac58eefa04a3b10ba2f786830a38082cbb",
      x"8746d5e986a4f8e3cbaaed2b163913ede3247c95b32a8cc9d61997146e87d390",
      x"dcd6cac8cccbe1ce2bf8220780f9ee7f130804a76579afc64752d07c96cc606e",
      x"af2429342aa6b0dda693954faf0ef433aeaf18870070be94ea22121e43fbab79",
      x"e9605658499ce0d7e93e6984d2b6dd07ff3a00b746a46aca7b79808dba038d87",
      x"995c1180b87d543a41ceab64ba3d0bd228ba7bdeb88826f125e3f1c9449b82d9",
      x"1fcf950d29c55114c8a9e8140a61d3cbd9eddd2f39af1bcfc8b93a3409660bb8",
      x"d9198cee5a69f5ed0992e6736e32f8714df37c0a6946d0d2fa798508f629fb97",
      x"e9018370ba3689f81a6277ab62aef142805d664d7116d3be9e23738eda071e00"
    ),
    (
      x"e1138eb2ea966f5e6b70e23366f188b38eadbaa60167645d90b91f466401bce3",
      x"40503e99d15f38f804cd865adcdae636775774c5d8e3312e72f0958b18c5ba40",
      x"f639b94f8ea287d7219311114d420f9dc28927a2341421dec221808fe0385aa1",
      x"b59d45fc8295911e08f2b342e6db70f21e9fa5978f303dce69ac2bbd1c0935ec",
      x"cfb9a9b9060823e0805157b3e583ddf3cad25db8b9446b43eb92bb816a52c400",
      x"98ae99c6eee1928d0dca6116d830877b201f214b47847d21c0d1642a33de4df0",
      x"d653aafdb5122e4681b2173fa33397411df9ce7e494dfc2b93f70a47072dcbe0",
      x"5ca513830a22b4df793ccd25b2e2c49b04518c3bbe83216fbbc09d0bb13d8bd9",
      x"726875354d6ef18907a1bbb8302edd634d586d60a726455790e47149659d23a0",
      x"2a87bdd67e3103009e627e3ce5abd145a4c78e173b90463c81cae5c49edbdb36",
      x"23018fb10447731ce30bde97116e3d36a4a8925a882584d9558a97d1cc2d6b37",
      x"d55d0579dd422fed32286d9ffa850487330a30f41a435a1a9d68bfa741743fdd",
      x"916cec394440c92eed4aaf318a9df4812b479059d0d8b57f007323e26ea16def",
      x"a7ac16bf982904c75ea36200ac919577fe8b5b2b5cc89590396ee94763ff74cc",
      x"72688914520fc92a7699cb9f35c115ef882812d4fc66bf2827e2182b8ed19b8c",
      x"28d5a524bb9ded89273a56348b532904fc0708f5d885c984a1d79bdc8cba6e6c",
      x"be821ab3db8701632533f87518a0dec8be988c5bc7476fece8909bcdaeea3c34",
      x"4cb132f3849b03e5474f6ad5d1dc936354d78fbb4fcbfa35d1338ec7d854acff",
      x"3a8bfedc9e67a5f65916a895cf5ca6973526cdf53aed19cd21d0ffdf3bd8d562",
      x"d2b9479d8f31d66ca63ca60c9f9eafdaac304f620e5be919c75c1854690f6943",
      x"87b12cf10d6f8d18cd8b656bff3967c6d11e68d1b1092e074bb26b8c1467f0a0",
      x"881648091e5a083194866ec24a8520aac71bfbffc94e5f2f90d54d3e705d0845",
      x"10410f35644d760abc28c890456de0688ab4dd374c41fbef4e729c0f6091dd8d",
      x"5696eb28647b95ed249455be27572d3e722f94877957259c75681b64ab8f05bc",
      x"14b9cbd2016ad616978cdc3286424412de0c17f4caa0fa72d0de15d84ce2b10d",
      x"9e42b84541d7403ab1d856fa2cf8dfd822387a2220da88d9ba8ccbbb0a03fd51",
      x"996f2daabb3c6efbcb3f5694d5d7b1cd2aaa31c24381b504419f1ebd484c90be",
      x"a765ece560def5c0318e3251fdf296d7881777c75c844079223b19b5912b996c",
      x"4ebcb6cd98a1a47d2a3e3c9d7c7abdcd861bff7f8b4c74d744589f0eb42439e5",
      x"3bea70a22cfc693698ef49ea39ab285caf6870c755d5cb79d93b11e1adc8ceaf"
    ),
    (
      x"411b173d4a8851e049f4b7030f12be5eeb607e44037737ce3d3452d228c7cd92",
      x"eb13fb980d99435c2b11fde6b723a98f8f208bd84714e723b3024d33050c2b72",
      x"6eaf916abdfd90514805fffe0b23b82712b902c5cc935feeb085923def23a537",
      x"c4cc685056b132b9f267d37739713329d22466f106e889062d7ee286135162b7",
      x"93ae6b79ba5218b313801942fb9173aa63b277198b3a180fbba4dce7eda465d5",
      x"3543ed787a30056c9b933b99f3b18a912838b78a474c65b9e13c3917ff6d54d1",
      x"366bb6d42de73674fed0c228c2cfed9c40f10cb24efe7e25bbaba2a3910017f9",
      x"75e8e4503b278698040262c87ca68623e1dbc267301437dff59948e98f5b61b0",
      x"d44c46838e1606d4968756ba7bfa5bb3ff8842f3b55024a401bb4cdaa7e779cb",
      x"c08f888423ff9a6ab0ab19b869a3c579f30db220b84125e506d88412a1cf8ca3",
      x"a662476019ccdb31629971112c772c633d72a776ebbd67db9c77d466f3551e67",
      x"f3612c52b620c2a639f2fc119e82d87b8916ed2a9958cf932a87705c616360e9",
      x"1a45eff2f7555d61750b38e473f4edd4e852915573a136ab4f0b740d2c1047cc",
      x"f2bf566002a3d6375b4e674369ea2825a9b82ad7ebfd79e3f7bfe9845e0d99ad",
      x"7abac39df41637ee0552cae72a12c5ecaa07e66fd9542b9683e8246472f6b0dd",
      x"ceb5f1ffd94bf170694c15b17d66e3a0558d645a530bc23f07a2ee6a7ad518aa",
      x"b8d77d4da32deeaf29a070dd6334f28d17454f59fce8f9866fd1c172f828cfc2",
      x"55b1e1d4bd86072d89edaa4c7b2cf8fd17ae6d23ebb7e968f6695ce072aea804",
      x"7f00aa2539ab7992707f079b8f463aad9e6fcd42708f10bdf54af2584d6464d1",
      x"7d4e88846de23434439f30ccfc00d3cfb749e7ac854d13f7a93624e4e2228751",
      x"57cea68fa231799f91215d4ce74afa9d40ec2bbc30ca433f501443b37e042473",
      x"3ce0d306d916f87dbb650383a11061cc20745c106b252123e8109936fa6b3f48",
      x"1bc8134571fb86aac8162d69cdbaf00ee923cc27b74452979a5933d9f2c8759d",
      x"5df09c459e399cd5d673609f9e3cda8c0838f3aa9eb82706ed623eb641335ffc",
      x"8c2282a25fb4c052da7c96b5adf44f1252d6fe2ef1decaa3b08549d506f467a5",
      x"4b55a9dda60ea6bbda78a2a102746e235d61e24b047637bf89fbde58f2064a2b",
      x"7709c43d79acec92da40595c1840c32d1554d93b3d94c96340896031feef3c53",
      x"4ccb94b1fda6ee9e0c68b1aa70787a5a703e3845277d466918c4444f83b4e576",
      x"d0a15caee96f5086cc7efc11df475f0045c3cd72335f63379849a1b94868b927",
      x"0476a715603de1b4620726b6f5ad2a84c6523158e9f9fb0f2781de9af0ac2a81"
    ),
    (
      x"9867c0c98620e604bfa5d3a9f4929890c8d62b49289000f64f92297688e1c371",
      x"87e1ef22e1c1c3255608f081f1dda28c2bcad8c331010bcc08b81961167ad999",
      x"9802c5e924fa5d81752eec9149e3ef65292983494938ca6dca041fcfe5ada6f9",
      x"c53c02add310756b1c749540e8b30b651d492c4ade45f7d5c851b7d7de75907b",
      x"863ff97904af9018e0e1516a098b3808d7dc072282d3a57dff1bce6d769ea851",
      x"d98d5b645f3171d91aec4fd34c528de03ba151e3057a3b1252d0cefd5dc3ed92",
      x"937dde27b21b6b560cceb30e371e4835d00bbede8443cefda4308743e6166db9",
      x"295b3d370711b4bc1bc11af86dc1f154b7d8ce6ae1743d622771f3f7f53ac41e",
      x"f88937eae892ba8e8c31e61dbd2fc2570f9cd13051a5f3794932dc9eef9fdb76",
      x"1d4055e0b3e49de384d0dd7be714c839c6cc7812d152ada8bdaff7e45d7a9da2",
      x"72e2bad07412c1daf5c79a5dcd72be1b82a5d1725684342d503c829485958f38",
      x"ae7de21343917a884399c30d0a82e8654aa2e524f250b6d56db49d9eb76efd23",
      x"55fe29838b437dce0602cedbb243d40ffaad95e9475835f3b7e5ae83e2e0d307",
      x"b21c22b2a782d32ae2c7835b8fd068b2b497671de028ea0bee03f58bbf637d26",
      x"5272e1d8da40ea871f8cf9d37298c3b48a9e1b61d9b97081bc9fa33a4cbac554",
      x"bb9de74faf2f4b059905764cb9137689f97498022e726c5cf37cefb8b4b38392",
      x"a064659e05ca08f65a24a9727ad4110ef3a1c421c5d178a6abb7c60234966e6f",
      x"c4c00ca6ea205a0a167164280b7e18c022c2208cd0758f1ad94b56d23b30bf0d",
      x"4326ae9541374b2c1de741e633bf7a3ad5dc8de2bd86d1a96d30218484d36129",
      x"0518a65424a509c83821671e8b85b237da9a2cd133e9f881f60693689aed8085",
      x"cc9af007fff85426234e4c6b620b31ea133fd7370db2f98f117f7c5ebf7139c1",
      x"ae6a3ba0225ba7bde9e6f5d241d207149820feefbf84e560fdbffb63d1ae8a5d",
      x"598e3e2115be877e652eb69076a3f6a1204c4b25f30421c118827f696e4851ed",
      x"c355574197c78ea1b10acbd7bbaedab45ddd4b5e8515567aa6690c95fb466103",
      x"8b1d30d750b57437758956e13ca000cbc80c2c66f0e2685f06e69c546d15e13a",
      x"0595bfdc15973e2774257be154396f2e358a3648e33636af28e43ce3c16aa2eb",
      x"0f4d5ff6383867eac4c55b080fc52e21cbf86acd7eea52691512ad5fcfadd5d7",
      x"eff9d9f2ee780ee6bf001792a95e36c56b1ddec9a50c78caa650730ae1fb75a9",
      x"968f0cc67c27fa4e74f766d591f4eafd02d8ed647eb4386c157a10863e11a174",
      x"0e6d77b450cf4ccd98bf42ea374c464ae25d7eb1674efd77a8d325e89bb3b478"
    ),
    (
      x"549ef93e607b2f99f35865a3d02d1725a53f458d78f7c364b105af961f117ccb",
      x"d136bdf4d10333dc42d4a1f443352dba4dc7eeb090dc13b719cd439519a2accc",
      x"2f1e6befc473e5a56c4982c9311748f6ffdeeaa4f177763d7087c2269a289795",
      x"b034a326bf51fccaf546211e6044c9eb9c2827611342deb96783d7aba7869cb6",
      x"b37ce167090ae40cfb5dab6b2e82fa8637412d38c524afc7fa985e3d826987ec",
      x"9ddfe7c57e9a32160d8033aab28c5c84e0b57a6c121f24a37fe84c5c6ca09c0c",
      x"4df4bb8c5281d3232f61a83052080cda37aedcb557f3533caa91cdb4d92fe483",
      x"dd7ba70653ecc48a3a860c28d83d22d1647e28de337195f887557e55e4bc3adb",
      x"232c77125fb9c56ead85b3125f7255585e9e0744dc492169764c664f349aaf39",
      x"e28accd268b5c25b55b25aee60562df675081594b9a1966e6f899fd1cf13660d",
      x"e219c6283156cef432e29cfae5ddb0b285dd0cb905737e7a2ea5a6d664018f45",
      x"ed27122811e97e72fa864d22488d25779053326bdbbcc5cfdaa631bbcdb87dc9",
      x"0f35df7ce62184ca186ad3f93c04659574ec622c6716884c479d462d5fbc3064",
      x"bdf6a16ae19ece6d25c0af41c5bbc21a738196d79371884ab2aae97de9210b58",
      x"aea12964a77227b4b3f6c3a1cfbf2716d667a715e598db8c2f645b797a6d5921",
      x"5bdae0ebb915af48283a33be1cdf94975acbc43ce8b588b2ad6170e7fbb7168f",
      x"3167fd289f818179c07f711f5e9bb4029ce23c693bf92db34e282857cabd04e5",
      x"fe86fbcc4588b46c4920c0f7e7477b5492e7b02685d277fc8399370f54feafae",
      x"063e29876c81e3928b187c1493c67ae9a50381b3c639b05a9a693a8266680ce3",
      x"1891bb10f1a429b64d1f8753a60b3b1b0a17dc0370e2fa09e041c71a4fbf289b",
      x"33991510254389596e52fa4dcebfb918d3deccbb9535c2a284d9bc11252e9ed2",
      x"61aa4e9c8f80dfa61efbaa1fef38530c08eb6fc8e315b96c80d93f3b7b8290a0",
      x"784cd1de32d1558a77c28071f3f2ed8a764ee6ad407206f79c51853570bdcc33",
      x"440a711f8f7eca89bbaa45bee40d85888cc4b197eadf772586b6049db2443e0d",
      x"9256c3d015f52f580d1fe140647eb107f8581f21fe5e326538346788dc9ac38f",
      x"164ecf9e3a0b43c4487b404d6b82d200cc6a1a68a4e7400c83ff3b7bccfc3016",
      x"2a89ac28569c5ef44982e9fe7dfeb4957ccffea4d3cde8a0c7c9dd31358232d5",
      x"dbb80794d1a388e78655424928e3a6dc305fa1fcd57b999d151eaa8d5871399c",
      x"015b6a0e6fd637692ceca96b0cc07379ef2836d89eb488b6cdb8755921138a61",
      x"d68ac287541ba5f0573d50fbd9aa59a70dba1dbd002ffd1a197f2cf7af511056"
    ),
    (
      x"4e263a0b8c3fca31195614271971228dfbad793515cf1d9efa9e8ddf8d08902b",
      x"81d2965ac967efce4207419a575209c41ea3bddce6533270bc281ebc31b0eb21",
      x"ee7b6a6ade8618f940b5a47bc3ad4b390ea51f50794ad3b3b2e9888f450dcd34",
      x"55eb4200036b8fac1dc7054361e4343fcea322b1fc7e604f7f48384377bf2a6e",
      x"e3a399bc409a3cf5d2f89d5668b17543e05378cb0904d295c6a27d49b97cb883",
      x"3d8db47bc828276d7a6e51c03236ea2c19762b3f7261333164402b7b515456c0",
      x"7fb4e0986f743dcac38b7abcd5364a6954ad21619c489776db653ab158f2be8c",
      x"8cabd5d97bc407eb06d3a31cce64891bc01cae3a6d9dc34f4ddce5e943c686cf",
      x"591980c33754015484c980f099d5039188d0a1e73c8ea5940d863e2c0353cb3d",
      x"aac62836cb79ba905193b66d5b82c00b910cf90b59f17efe18ffce5545aa76d2",
      x"b8270e4271a4555b8086ed60e642d696089e1cf5a48f2d8c65fa25400027bd7c",
      x"07c61eba1043ebc54d122d115ea1945e4c06b31f2934363fbce44d85ebf30ab2",
      x"a044b06f63123999109379444b22a1b1224a79878df3739b2b99e69945c5c127",
      x"0614091ff2a504ce70fed88d7820fcc5ce2fd61c95204fbcfe6045d2e35cf472",
      x"5e8014f30a789266517d96da414a529798087931e6bdf173f8e455f9c71d97f2",
      x"ba0ae1d11c496bb3a802635daaa831828e7607002b4790bb2536b36bb7e109e4",
      x"d67389f87ed74cc50e901eda4a7e21d7ee1b4f7c7fc0d0c7598e33b58e4519e7",
      x"4b06737ff6004ad8f20ee4daf48cf18b496df08f7426395abd249cf112926123",
      x"7aed971044a13ae511d1075431ce91162399c64faf9a9d994b6c57936f4969e6",
      x"9c6dc1df7a4be12837e4361a5f71ad892ce4c63a9e73d2f32d10ff9dcff52ec1",
      x"52800faaf5435b0ed706e20f8a42ee3bd769060324f2900e0875361aebf30bc9",
      x"3df6b7fe7d12284124f423db7ce4487eba8b69dc42e3b0230345c152bebafb10",
      x"d3ec1a6dcebc16e070df759cc930a34137ed51feaa3735db155bc03b8e4547eb",
      x"65ce1dae730d0183cc323a7f857747b99cd2307af75e0d7df1b0240e2c9d5868",
      x"404edee71bcb558e43b7cdcc927a85d65ccbe8a7702bd029f1974dd29235b5c7",
      x"950b5b0c8e2570136853e60483543b648baf4e3cb87bf1989e2698da5aac0b95",
      x"6b5fb12f948fa93f82430fc5091155a0b52031029eb1e20446e1bc992a145a15",
      x"8623b283c9660dbeab79b1bdd6b571de80101756891d053ccbbd02127a89c121",
      x"c0d9e61d5c84824d41d929f10d998655026d7ded8d87a53913650116fe5bc17a",
      x"aa0cc25fa03a1d0d336ec17eff742927596950d3c969890b51a83dc5c00444c8"
    ),
    (
      x"bd5c366a377e5195fb47400a29e7e29207ef3289e8ad293c80910e7fe8aed325",
      x"1683fba6a27c66f6bb10e8eaed15c4f4eb4850604616974a29b62b80f7fb0421",
      x"1168b3284010f4d2c341a329d147e1720bfdad60a272903a0bbb7f3e3b37b45f",
      x"e54b570e26b42f67c1bf6a02eea3bd0a246bb31c19068bddf436d746e7cf7856",
      x"3ee9f6837fdb66949949b4670a0594126e80eaa7f8b3b70fe3ace8d4ae8d3a23",
      x"2c9f48728dc0d65ebfd8c27a02806505adf3dfa44f197172ee428be26be15c1e",
      x"bbe60442ba6d6a67cd37505efd28ec7136fd37534de1934900c332f729f0e944",
      x"cf139cdf8f88c660741d1c4eb96d3aa8e25fcec1ce0a8f29022401fc04ae6c3c",
      x"9aab8d8af402841872b7f6860ed5f8321c5a459f9a46208b708cd233036f879e",
      x"0bab0a542716ef5e15b107a172c20d9b19fbe65316ca94888ba882492ef28abd",
      x"656b273896450b130cecd61060cd11bc68b641794044075a9e7e5ad6e64bb791",
      x"5fc4c257d8a2841015bc1ad809821efb1f6011922d238d5b64b3e903db3f605d",
      x"bcc5099d31d8b7205b987d49a6870d4f51c4b744ea221328e71334a8ec3841d0",
      x"6157b2cf9814ab408006468c547886f7c83a54ad6d3e25f2dd98261959af587b",
      x"3d796b8d8b8baf8c47e187d03da28cff6af23d908bd6c93ef50e43b074e9c9e8",
      x"cbf8e221ac1d59566507b4c5f115a6316f7c80e845c5bf6a55df9ab9e8472096",
      x"a6689b85ea28cf025d35b7fc78cd12acec21e9fe972969d9b08632c72ef86f2d",
      x"dd880172f2b422db4f0fcf2d031f06f523df18f17d308e11978203d5dca97a89",
      x"d499c37c4ff122a081859fba003b03e938db4f0dafb27171967dc2a2bcb8810c",
      x"453a110c4e4c88b9f416ae5f4c1f2ab46f4690772ea7e270308be6124abfa7ea",
      x"23685639903953cdd0ee1fd8bc570b2289643b25185fe5bb98268c2d5ddb15da",
      x"f79b61989744100ac53259a2a88255249bbab668cf79e4f9ee74df63681507e6",
      x"683763758876f4a23da6c13da6751ce5fa5bb5d37207c033f8af75fd34a8ea91",
      x"2c40128ee9f76426f8af52834c8f5adc141d833bdf513fc3e4e9f440e1656509",
      x"06c378bc9deeb5c9b313364b730a9babe79ddba81cf80db68a1b28c734b12931",
      x"9867d152276f7bfff0bb2b1ef557e2b5796c84c99df4202146fc57cc5c934bae",
      x"c1e674defc15c09833ae848f9ab59a94a29ef3e1b5d44d320dc30caff134e822",
      x"e51b9cc706d8a3d64a36b9644a58944847dfaafc20de1ed578c0b1389032873e",
      x"01c4b288e2d762f551e8815d74dca27d9e0ffd2f0f9ed3be465fdca0f5dd08bb",
      x"ae87aabb8eef08a7f2406beca094ace704730f936885294ec59559458a614376"
    ),
    (
      x"1ad1076f04ee9598f627e33e0b6fbd5ae0e876e837282b97c8c5de20660ca910",
      x"ffec92b956e6c972c575f3b0c2cd664dda6105c143d40d503f6ca98584d528fe",
      x"f5b1b6011fc1fd44cd00d41b3b05633a5128c503c44d39f205da83e50664cf84",
      x"95ef0289bf677c63c0661623a040b75550262749f705c3aa14361410acb80678",
      x"80fa4ab1a0fb3dea8699b77858e3d397960121273ca7389e1ae8ee82e3c8c51e",
      x"756819e2a9448131416a085ae82150a0d6424a5ce20ba74bd3d2c256b531c208",
      x"3e842459b77db57b10ca77dceeb4e9bc0d12266be166d0a34eb7fe3cb6fda6e9",
      x"1d2b2b7a4aafe77cc493834b4f42ffc2fc74b8576e0a74f1d3cbeb7b0bd449b2",
      x"103d5bcec2934c5a513fbd87ebc2967ec7ad0767671ac1e94a4d5bad45378556",
      x"f92f9199aeeeec0ed1917989277f23b0e23744670ba9ddfd3574207384909434",
      x"5f2f80b4fb3822f1d1e04b8650bf32faca2e14f6010899a34068aa1d3c723462",
      x"27bff025868bd5f3c0ca43f31317c05f69b5fb0b00771e083b0684f292d08953",
      x"4d3731c25ff54046a27abbedcce638a1965d054daa3c4ea3d3dbd5f645e38319",
      x"331c3028456722fc18fa97c80c3753c52fb08e0baddb04b16dca6a44cdf65bb9",
      x"ab3c6af78af3f84a2e089c293ceb449c47fdbb2d76969c022f1584c5517dd2e4",
      x"c40b8be6f732314aa01c8d1b17fbe2bf0bd9389c9b48e6986efc6108ca82edb9",
      x"c81c435bd885f4fbe88021619bb214673d67bae0a0c504687183fe210b0bff3d",
      x"6261304bae3730bf7105c586519c5b21bb39f99ebc2ff80cae7bdfc68132e2ca",
      x"8046a8a7e30729482118f1a62c9ccfec2b6568de8d47d4f27f9e55250715ad04",
      x"d71b18bde0165097f243890dc81e88e33ce4f7d0d764a4c58df5c943c78184c5",
      x"e70bd96c1e22bd652107ba39f9f69f06395b8b9b40baf91e6f96bb5bd786de5e",
      x"ca8e7ee4c4ebf2d0d0b065d21626ca5047865eb25bc88a35b8e0ec410c93dfaa",
      x"e9011f7eb426dbc06d2a8115bf3c5a4a76b338e12b6cc7373deb9e987b4095d3",
      x"826ecd1f29a67e5fb7f7a74f97fc4591d892830556c930ece11df0e1971ff2f4",
      x"88d209f3330dfa096e0357c6650a81c099b7432e98daa9e02461d9ad8c6dc915",
      x"14fd183c9bc7e37b186d8a148c858e2042a865599fbb09bd2b025ce4e46a3f42",
      x"bf7f4056340eb5d6ad3260f792bc1e6316c1745e9142fd2f11399567156850d2",
      x"e483fcad27569e9af50f92a0b5d7b425755d11171b3f3cdc78db1d848404673d",
      x"63608740187c1896f50ca4463cf5a2a6cad026fabb0c47cdae271b0faf10b081",
      x"0dd6543755b984b7cee9ea7896ff91b6fb9791ee7c0f90b4cf127c76d9f30e39"
    ),
    (
      x"197626ed705727a10e5c1f01471849402507ce5730a499f6e113ed264204c89e",
      x"28231875dc10f6afdb8314f125b533a2e9f461ae63cc3c4a72ea3d4c91e1bc0f",
      x"e6ec426ef78d1edfc8ba9ecee4b57a22437beb1c047c3bfeb1ffe12685ceb474",
      x"85b72653fdd2ca2f1ff4f005cae23df66ce3255f950be4a79af35d9756e760f6",
      x"65e9cb48b713da3bfc8d8cdb7bc943cbdce473d8e2b54d859be58ac00396ccf3",
      x"5ce02414561c7f15a61773faa62e490c226577056774a7f9b9a9a52757224f31",
      x"098d22fab6b754be8e581d9d20242964224e8ad90febe98b23e387f378d1b4e0",
      x"fb94937dba2470540dbb5839ed838acaeb6015481a1077ded63e9534be8785ef",
      x"480f7d0321e3c29a326beedebe9142602f207f4e140184e57be57cd83a1924ca",
      x"786ef53679396444598a94af3d1c5a976da745bb4985a42c1f5ec5276962d94e",
      x"554136f8824f2b385b5c79300b645b628b66dca117e58b18743e8860f2f27a5b",
      x"a09302c86da4a75a75899cee29aa9592f35125bba28ae8481fae7998be0ab6ce",
      x"0ec471ed7775580e73ef173afac026a49e098c65daf490524128da556e38cc3a",
      x"ab962999a9e342b004a9d5cd375d49b240e72e02ea592432bd392afb15beb652",
      x"e8f69621555cc2bb2c8548304ea9b85b3ef4700f77a0340962f4c5bd2c2b82d7",
      x"f09dc5f8be6ab7f0f96fd2fc58d7c8a31c778dcbbb87cc072113c91b7f221665",
      x"a24922c7f4c1f3834eed3b8f20492e39fd1e8f85e3db09fa38293d6f417632f2",
      x"0a9e3767b7ecdf734e8456a44786c5a481400e5dd7adb6fde88c82f42939bac7",
      x"f8b48309403fbd7b2977f50635a52776b36a581d2db628be93451ca4dbec5530",
      x"0dd243d8edc32eee8f31c86bbcd8bfc3938ae6f453974c0b47522d9731c21048",
      x"e9a1ac9d4272754ed43800d48db00c935697ba8a5081b3373677f736f22ff9f0",
      x"95d20acd240d998e692893a741d1da0785d14e583eb8eca994c33c5af408ffe3",
      x"e7f544f6c6177ff81c18397cfb6ca34a2f6071d888edf7a530ceef55da1f2ce1",
      x"8cf1349bf8c61788ac778551a13b8b6bff9553e2c388468eaf500e5995e979bc",
      x"ee5b397ee78db11c322cff39c4aafd5b23655a502df9148fb15b3c806a6ce411",
      x"4eca9a7f5784bea0f15214f3c84e36ff357f1daaae1debd9f59a7af88c5eaa31",
      x"6f05f90d6b9b928cf465e3c18f00e0db4fc1c1341d55eb826f4508ab1ba3ca34",
      x"5600755a6a27738d578f2729339fd9eba5239e8546e36b3f5d709bf7263c8ef4",
      x"3f653ecceb84b4170019ff00af486fc03f0978305114a9167f24d10ba47c8e5d",
      x"c24a2a347ebac48d038494b4209d93e9a31a08555ddfd6f9ce67313e932a28f7"
    ),
    (
      x"ef3f5c84484944bf12006ee1e78594297e5ac9286e3b1e0b6012fdf2d0f27dfa",
      x"1500c33877163490a87f006e1a3fa830f09d8aa720ad85176f82a01fd2480d6f",
      x"ff1cb9ad7e53f06fe100450dabb570c6bf974f6abbfaef0aa5d1b6b67a86ec21",
      x"7c2d5f91e4e1da50b2aa35eda64b1794b5a7eba125377d5a0362fbfca00aaa06",
      x"447012895333de2d8c12582e42cda3e87ed36be08283b91432e93ef2b569b776",
      x"027224b34f73f8766833c56cb1831b5c8da877ef3b0c7e7c3c40a512a4011546",
      x"51427b4ca253d739bd87e6b1daef29856badda8fb728f15a2846b7bfeec4f237",
      x"48544dde8745899a754798c46eecbe0266d8aa0f81a991d5fdb7b4d3f9800bd5",
      x"ba2dc42f993725c5bc6c9c30f2e1cabc95327dd6cc8643e75a4dfdedac3c417f",
      x"46042562cf227dc28aaf6ef162a98652b67c902c41235b44591793eb08ab8bb1",
      x"1dcaa1161394f7f5297a55754eb94cd35f87b3f5f60b5049ff39d727bec578c0",
      x"d15a8466d19d2916ada90df91fc4595793f9be00b869ba8b5bbc95b12195fe89",
      x"d7b3ca9fe6e48774baf210f2b19813c27ac7c0efdf9dc1013180798ace91c83e",
      x"01ccde44e9de3c269e7c9beb4a9988a88037b477ba3d576adb0140564b512c03",
      x"83e991d1ff4a21179930e29fbf1602a8b3964640ef2fa126db80d194dc8f0cdc",
      x"791f58bee890a9f79e7a581b96e429444c62d8ee99ce59c13ad622895993e036",
      x"a700cc53c30a4dd1e65af17d7fa6608013c25ef4082ddd60fcccffb1712ca712",
      x"6e38110fd6a3834cbbc0aea78a634938dec5223e55c8d7c73ceb61553e2457eb",
      x"dc31a4972e7066db3436c6caf79c176f714a2785b89290f2e860f5d628a6bec9",
      x"806350bffa27cb3d4d909dd9358862ab45aae78d6d45afcbd0cbe69ecac6c529",
      x"0a1e9243093e3dcd8c520c62d9e021a8a5f862f0d910c4c48ab5f42051a87276",
      x"0e35bbdd1c07fe182f0e9c2b09f50c0be0cc628dca1bfc700ec4d8537e2a2e56",
      x"6a95f1a785fef70b8b1eff5040ddd9195c856da6adcb84234671d719492b3588",
      x"5f1ef9c9bd08f5cde531d21239372644fefa575e86220a8edc88441271f69c2b",
      x"1bc949a54184a88aef899d2b094adb8f783e8a4ee1f4b13c8d7f2a0d1fc4d349",
      x"20ed383773a2acb96f47092fbb31968785e478054fdc20bb636b581dbf4b8a52",
      x"9422bd04cc032ea2999c63fc4caee2e473aadb57ae2e87e98c5dce713fa54f9b",
      x"bfef35fcbe4e324f81ea69b12e53db5dc01cc8097aaf74370dc311cdf6281e66",
      x"2180b6754b9a2b5944506b2c3d13a8a98c805461967cfb210c8f4b198077b1fb",
      x"d052715dacb3f9665c08d1429c799fe6c312fdf7b8d7d8329abd72df8f7c2b15"
    ),
    (
      x"a498b2c16eb7330a17c436ecdb292ab73ba3f10eb9c50c7f650bac86ed6165ae",
      x"19b6aeba4eda996f03aa2285cc0c6fc0adec522bb7921c849fb4e75123daf1a1",
      x"6bf1d5fafcdba9f4382f18a12969e0adf7d8987b35a361286eac79550d7c8622",
      x"c2bbc6caff1c19e27237dfdcc983bb84bd712be40c5b2c49f764aa4581aa7d46",
      x"d3ed75d2ffad3f653a8cb54435c2a64a0c3dd3116b447a46d0af5d1ee38f2e50",
      x"826134a4897287e0fe171f050ef989b95e842eddde26994c652c44700b540906",
      x"586ed564ed2190975c53fb772d4210929a316abc67f11639dd12c71c1cd834bf",
      x"6a3878d43885fc8608cb1b56583fb2fab095f8a607220d3f03b3e3f095a4ea7d",
      x"5071b2dc7e1b34dc9923fdc7e5bfa0733d24a33d69d4f907e229899dd78be3c8",
      x"26835c81f680596cf60c41917eb46065f74c65a0490f458794344ff2ff11e8c8",
      x"fa158014eb2703bb88cda4b403f6dd5a1ec388328722078e72d62807b3a750f6",
      x"01fde50a03cf52ec4598dbe833427ed0152b22b429a9e7e8537b80002e61d066",
      x"1e45e68fc9eec167178498f11bd83b1d6135ed497fc2cba124a6c3e033d8f6e5",
      x"629373deb0e4db3058dee13b6ca1da832a93475cdd3f4addeee1756219cf3aba",
      x"787beea9ac8b9ce646e7869fbe0caebed5df07f56c34a58aafbbafa7634d255a",
      x"ef8226ab28f9063c94202620657c8dffd0206358f8945be1530e263eb8c64293",
      x"e6f4709673870a8abbf2972da27926fcf2b48a35799e97fd5563fa51fe385624",
      x"cec6a8ecdace02f9c81429f4bb28acb2c42fb0ce8d1e56c31419748e142061e0",
      x"de7a064d6c66b4e297615528fec57834a1058f6a51f08bc12fce437c28adf035",
      x"c80719016076eb860d3be2627f3c9d12f6ad393ce3cba22f5d3211d2b92afef3",
      x"4af74766af94f546968cf787004fa98c37c89b737ad57325ccb62f9d28df8179",
      x"35aac8745a7f5744583ec3d48a2425469f3295eef9a07e052671fe10117531bf",
      x"d549c94529924046ef6f159cc17647f7847e2ade3ca176b2c11878fbb26600f7",
      x"c72a3ca1c459a3413c8c503c00fdeb4bb60dc3567cc4812e0f5ed880ccab657f",
      x"2869a4221dc3001e3da87247257c8d46d11b9acdf324929a00079898089bf041",
      x"dc0e58b8c8646c19130711d26e361e2ba6e21709da29a57b7820ade5bc80bd5a",
      x"380cad4b0a4f441a4c10eb7ee38f41919ddae505a577767e483454eba3dcedf9",
      x"6fdb3e9580560f4234a51cbd0566eed3179f0a06eedfc651e0bf2ea0106affcb",
      x"966181927981e8dc62a0be7fd2ca9030409ce5b9c064fe6750a6f3a1e9b846f2",
      x"f367dc10de1effeb79d3bdf668f702bd94882415aa2982b0ee8de2c3d9325e43"
    ),
    (
      x"4ee973412ff211c2b5c6e6decc7e04b397ec1e92acdf4b98fe1391414eac77ef",
      x"2d52980aa56549a164100edca4c749ab6565ee3ccc17e63dbe045d3a2f0e3fd6",
      x"bd552c3e23dd817b44c9e7043077e6045ccff4fc2993fc4427dbbd65cdece975",
      x"72c5a881546939ad692a02cec51c21cc9d5a4481929bae8a810197987b336e97",
      x"4bc7098bd65ca130d2c93af9043b4550f956b8d65957a3bf29f4870ace5876fd",
      x"898f6ed1be83df45a7a98d5b619ca0027600c0b366efadbd8737e9457cbd9f7c",
      x"220be7437c1d5f87c7c273df188140938a28ddba22d1985df79e28dca9bbe22f",
      x"ed32f6109b802d838b87500d11745672b9d7844ab29bac8deedbff4a5a193cd7",
      x"52f346b0d5771982994281dbb3c6f55e7c9f2745f5ba52511fa283cc4d6629d8",
      x"fb16e45a5ea499ef7f45f3b64f868f2268b49a40a88b7bf10f4039af4cdd1ac7",
      x"cbcd0fdd331354cbac81c243d5c2366ba63e67f2c45757ec2aac30c7b8959791",
      x"95acec902c96ec466c5f60c8078d89e69d31f2d41009141af09704e29ea5b914",
      x"d3d4b1efffc10817098eaa2ed027fa5d2a61cbea8daaef65a8ca2c37e8130d33",
      x"4da570a4ac2ed6808563daad39d930053944550efc623f43b412805c7c7b2c24",
      x"59f987423098ee46b3e29c20dbe15c93249d1e9163d125d4b3046caaa4d99f0d",
      x"33921648e9f631a22007588f18f0174818add123cc832f341b7c368a0c28660b",
      x"95d377eab40824b3266e8179708d4016c3175d25a5c8cf7411c7c7d0b86ceecf",
      x"fdd12ae8c8ea8f663d279757ddded08a939bf372d854e306bedac781c72625fb",
      x"77af5a77832de30d548eb30a7c93dee3b41aa137b3449eb9e45dea173eca2f9d",
      x"d4a7c74c25f5259d496c20eb32d63be283e09a89f2537b0638fb2c2eafacaa63",
      x"9fef7e042f562d6bfb063630330fdbbda08cc31c6279482380c5cc94df0999af",
      x"48c0b05cff5206ea9f9ef48e2118e66b85b415e917ed9c0e5ebc479226e60a57",
      x"709098b4a18a6509928c88a0f661353d258bf98160231021528a332f0c2f1608",
      x"287b950c20655a2d442a51257ca49ea97bf766b7bb0b691ae598daa4b7ec0bd5",
      x"07e9af2133ed5d5838c43e0f1e99c7373a6e0fb1589796cb958876d080aed884",
      x"b73e079f1995d082b8f58b4597b5d4803fa255df97f812d942949024f44120cf",
      x"0d79ad4a01081863fd96c64727b4e0532d4c0e7bc320d5c76e6d703505eb0fed",
      x"709e0de3f3c17ee8d7d251ee3fef30eb259f44337746fef16a392696dfec5f3f",
      x"ebcd224773d070711aac8506a437120a552b78161bffdc85998ef4d7d39b6a46",
      x"b955d68a80ef79e14dea573678d5df139c4cda897a096c8b7b69640fdb75ae24"
    ),
    (
      x"feea46b72abbf8af9c752c2c1021fcc5cce66c09ed2d1478c422f1d8600e3bc0",
      x"5483261159f55d69b27522c5ae4ec8b420d04408bd93c4229cd9c7647c4a4974",
      x"6f8c6d8f9ba70f81cb1b756a0750ab52e61247d61b5d244e374945a480e0384a",
      x"ca4ce532c1a0787d1733150d03ae14411f41e9ac2d59b6a6a5b64c01c4dd02e1",
      x"5986033a01fc9d5eb0e8fc35408519af94fb46cccc01d7b5eea080603f19a206",
      x"be61a03b0568e536bed7b99d5046ffc2932a680fbb42e7f655795cd4160364aa",
      x"dfc6859208b4a99475ff9e3ad400f19dd309f146a3c9b8ae984ac51f4c6149f7",
      x"e9caa4ac482198c81823f5ecd4a93eaa720d42c08512a5ec4e80148ef6dd7e8d",
      x"11ec37ca125fc8a8d0edc91899f807c58d6ba0cd963ac9e323faa2d4dd1e4edd",
      x"6bffc7d68176706a4e21f7599dc4a2a54c1009656f839683c96566f85dadd5d5",
      x"33efe7be0f15d56aff194d25ecb7f7f5b61698f5b9927b36d75a1a4d72d4fc2b",
      x"8a4935d616005bce4de9fdc49f3a327bffd885b16a4dc97dd26abf0b55914ada",
      x"78bd2133ed54ebb11ba7fb14e00aa72bfc1b27de9c21e7eb76cdbe8d9bb7172e",
      x"5aa370eedbe615b7083455af3a2487944ff5516e86149ab949a3374773654301",
      x"7f1faa672367ad87e173307648d4e88e6474afbd735ec43dcaba23334c590bf2",
      x"70f1b584f6dc23994ab5a62b734563c791963087573b795954db14e8dfd2ec54",
      x"03f785a85e2075dc243ead24ffb017027215247469e5337bbbf127fe85c15d91",
      x"feb79d5a62092e76cbb73475392ffac2605970d09ebbf7b136205ad00781fcf2",
      x"64364a1e7785a8c558a9a59d089eb53c083ac29d3204d94e637fdc690b331bf1",
      x"9b23c7d6da5c92aeded6dfdaa760a66e32f6f2f35218866cb0707d9caf0dba69",
      x"ce2928433ae27f29524405366cf13203c0baeee81c399052b5cdb24ac0476af4",
      x"714876830a76132cbbc35b02535cd510a9aaa222702be4cae81d339c902e97b5",
      x"006d11a01f8aec2ab59f5840a591a55f4a1338b6e4144132959b5ed6880f7275",
      x"e3bbafe858fb4e9c8c4d9d008308a826f778e230ae7fa88c7b70e42a498ee274",
      x"4ec1aaa101336fa4480b7ad1f265b0183ad5e7cffac25686c08cb95b56cd9d0a",
      x"81370687f65ce4a8ff8e87d3b21e1fa705138ca32bbc7ba858da2002d9537654",
      x"b0b2b203d6d5dcf556a3f62665d277fcc1e6c5297aa949d51d4943fcb2e2fc9e",
      x"72ca024db7613cc231eb1e632f04179c745d59e400e0350039d9335f3b541973",
      x"2af99fad6a0f7c34abf90583b432280670dc99bd2d8a9fd2b9c1028048a95902",
      x"11baed4f848e08459b3f5da01d05fd95a3937bfa450d4bfd77d1139a0e57c866"
    ),
    (
      x"89b1bd1f772b7039110af5d14e110a620befe3169d17f391a44f84a78e566733",
      x"2cd9721759cb4dee469c3e9d6a00efc5578a48179ecff075a836a027e9297d15",
      x"25e5bbda612b188ec8649de6340de648338a910be07720841441dcec3731d9d5",
      x"93f97e65d228ed806267723462b735eccfcbd531e3b54585a92fd61d84ead65b",
      x"2d90b34ec6b891fea85bf37cc449db964318c352d114211497ea9cd4b24f7812",
      x"adabcfd3a44239d83081330cda7b8e00f98f530df9f48f10b1d0c576bbb7d770",
      x"255f2e1aa80376047599b75ab2830862590dacd1c84b2985d15dabaa8c658ca8",
      x"a61082c83b7d61f2eb35279e2b4095372c3c74af806a2e5e06c4d61ae1f6c60a",
      x"5ae2b3a472fb5dbb0df332075f85fd680afb7a3d82fb72bf1acbbae949f00ae9",
      x"181d5e9407be03eea95fd05a9d3e2a387271c7f5c1408c34f19d7404caa95df4",
      x"1b9120eac95b4d3f3a11f36b5b63c786b28c3b1d6e0429d7d47a2f0a9c0f6444",
      x"9236a41f85a27a60180eedafebf707df18c004b13cffe0296308d2280fd66ed8",
      x"1389ae10ae3c59d57f9a2e66212b79bd5e7720fdd764d9ed2c1b0cd49061e15e",
      x"ef0839bcf02003ea8a31605aaa924888de5093fbbd8daaf76f306cee9b4c68f4",
      x"c0dab8cc68d3dfe7fb009028138c767ec42a5bcc7f2091c321c6a6cb641f4576",
      x"f700932947ee6fc1d12d9dec22cfbc35f80beca86770f54906133b04534ebacc",
      x"7749a16eee0841244b16871249fdc9ac944f0fab9c1ceb550eaca5fa88d58338",
      x"e7a74566d0dd9282255b15da8e46065ffff821e1441579ccdd9cefe117728e42",
      x"4b08e1d124b28592548a1cca3e8185be00fa80ade4177e018a4117a35fbf73e8",
      x"4318ae117a076e1749af9660271b9ed8eaf4dcd0c6726e61ca83b9089e60dfda",
      x"a2ce183d52e1e1713b9e9f18c3d33d2a00e27626d9d255c3fcc7e9d62c1292fb",
      x"7c968d8b870bbba00e1ebac84dc61ba9a7111419b034e4e3f571a9cc1a3a5a9a",
      x"57533577beaa29df53b2aa95a009f1d0f78cf8a4de1ef7fd25a5be0c929babbe",
      x"99e5bb2c2749db6315dc948961509b29c2dc0f441340a3a9907d4c3383868bae",
      x"ad51c06dc76ba052a382fd85c8318569c6230089848b3a6ba4e333cb60e159c1",
      x"431d111c99444693840477c0416528cca05a7949616a7a2fc675b3ed416628de",
      x"5885b6b688cd68004c613837474a9bf11a4f181d894e5c485fab767ee1c813f1",
      x"4d75e81e1807ee045b2a85c418b61471de03df5f6880e9d71cef9bef1b9cbb3d",
      x"a2ed8e97d59a38f34614982f4206b8c7e1901d71bad559ea471fc41bd6ef7855",
      x"bb68fcff6533aaa3fc4e6c2779c7a3fd9ed8970668add65cb2c0a4d7268a7a26"
    ),
    (
      x"649f799a7619992bb792a576e9be6939a6cf972ee52f4e56a23abb38dd23aaf1",
      x"3da464e5acf90864b3707aa71603d4a507989a3e59c42d4240e85581ee509644",
      x"3980647231c9aa98e1273f49f10218ae216d7bc428b31a1624fb1563c133bbd4",
      x"dc04ab86788eca13088b381382e26e218cdce659401d21e4c40dc3563b4d740f",
      x"656e39ce916811844672cd4777229f4f791563d631d81d143254bc18da10f7d4",
      x"d21c638115d4dd6ef3e6a4a6b6567d6f4c3b041fb3ce5b427fea5c795f54c6b4",
      x"b7eff51d167ae4a2c82bc59323d17245d824abac4f40d4612ed2f04f80469507",
      x"a6fb29ca8281a5cf94f0831cfb6a1691d2900b4b43ea19aee2fec86bf0f57fb9",
      x"fc3e4f994355cd9977550d5738af8e042ceefd96ffd25c27ec0dd5a205e440e0",
      x"c819758edeb0b90883893f7f09cfbed23b47a6b2465d22cc51cab67e083f665b",
      x"246e252d13b009785050ebfc82e93432e43cee01efeda59c51a604c4dbf626c3",
      x"2aa728a5d2732c0a027bae673fe71202d65be141e165965fc8d7ae3760d37e31",
      x"da2065cb487ecf0d081ae05385a0539b69da704b1ec0b9f3a71b802d18a39fea",
      x"5a8ba7fbda57f35ed83407850a2e8c2ab137a6dd6c5f605b18462ca2e5d5c6ab",
      x"e0ffb68cf7a7c6611ed577c631afcdea61f0a4789137c5189c2d25d4b5d64821",
      x"8488cdfe2a9cf7f2a1d188ca44a6d19c597b22e350704617c54da9c02a7a9a8d",
      x"b800184c65d702a2ffcefe3ef6c0739beef2e0843acb4cca59039117e2bc9b7d",
      x"e267dae2b87f127a0b73c69d93301532c9067beaff5a629a302000a63bb4f672",
      x"3c27e4c5a35d013b8b0e390520c3ff8be7f9f765e2156d89bc8284602e5d49a8",
      x"85c95c663fa6b7ceeeb5d01469e3f3577e4874bce366dc95fd73edadd6305c46",
      x"64e7e4124b5774017b6c434faa37b3fd1a8393b384a4465e8da16e17806c1e54",
      x"e84bd4e2211ef2788e50fe65c8b34e69ad755be5a757983cb2d9d8ba7727e7b6",
      x"f15cd98ed61617c5c5ea9ba8f97443541a7222117ef2fab781ab5fd0d585ff52",
      x"243a809b83385172aa5deefc5ddafe799e75a9597dc641b0a5833e71fc511988",
      x"d8acc56227883e9e6c50004f19cb8118d3c6fbebdaadec61d504ce7e531b5d86",
      x"3e9f779f5a3eabfe4f9ec9842a2528154590631bca10bc694f26576dbbbec048",
      x"d0688ce8cbec353c9b29fcbb18521d53f71215e2eacc4ca1901d6a6919d7133d",
      x"ad631276b516dcadaed0f37e02ab76a2b6a44d167bc6efac4a552a66662cadbb",
      x"d636e76711d9b107e74c40ac27e798b687ea61def0e74d77d4050011c08b0e25",
      x"ec2df0cf50d1ca0129d1c2649da339c01e97878c0fd621aefe0e5a3aa58ec5b7"
    ),
    (
      x"8eff67c59827111f514c2e1c27b264c0756a9932f299028c9dac54e698cdddd7",
      x"542ae71ae7495cbafa171b0d8e34e02053d40e8b90cc51eafeb752bc91d67d3c",
      x"7151f9c36a49c91dda14cfdd304d208c8dfa79ed12b9703cb186126c9c88ab71",
      x"5cd002f7645ce2846e2f5c0cf1dada1224ced55eaf9bb5e3ffdf74fa14b9a9e1",
      x"6568fc04e44e0a079f923f69586d690a14870f7611f6a4c4bcfad49cead45186",
      x"5a87d4b122353914a94d51a52ab3ac982409c9793a5f0a380c72a9acd635850d",
      x"f70b0771f4edd5e430365195c0c32c96e4cf38f1e20c465c2e869a95ea1440b1",
      x"eedece9a6cc31fd6ad89640ccb4d32e7c8178e15b845ba8114eee5a7d79a51f9",
      x"fcddf485ce3e6266a44f56da255cb8ea8866abc7ac73fb1ca05274e9b2138a60",
      x"cff8c6d26572a9401270eea1731e8d57cecee0de49a8f441534f4fb5f7650122",
      x"1416ef0769903bd48507189de008aa5bd4568a902441c57ab389c8749e45567c",
      x"46e576dc38e3b51228627d60e6686fd45570fd4724ed05f1e7cf88b703bf66b1",
      x"780d7db52c1d7af9590765a50f85774a569a2b9b9dac03ae9733cc3d6bad50fa",
      x"d45327cf75cd7bbb8304e8f9c10bdc3c16ce1d6e53c70c68392e3a2c680844cb",
      x"c7a7db553578018a62198937f298800b3de6c5d70f5a2a1681670425210a3d4b",
      x"a2ef21ab66410db9582aa5dcf7eda231f2b37c7bed8bf32e9549a7118912da9c",
      x"a7e054d63aac53605824042cacc75d957e5915b30993e146bb24f6fb33a4f8b5",
      x"ff5b9a50c3e53f206729be3881e0c77ce1456e8f3863f78b8b96c10c9f87ac0e",
      x"6c4c6e21f3e62bc79862325d1620703a9d3d163bf0c17a9bfd4e15299ac10cdf",
      x"bfea6e2be3049e78ff8e7067e7482312fca4c6eea67276018244247aca1e7b3b",
      x"48caab2ac626c6230a81165d18e6d261b212e72477807cf8db87888103559982",
      x"249329654dd959fb35a5c07791baf8d84a38d5721dfc1fb798dd580803f6cfc2",
      x"94175bbe87bf9597b023129014f1b9fdfdd228b8f9901e362176a9df7e53b2cb",
      x"8376db0a15c56ac0213867bf5da6fe8070c92f3b2753db28a1493244dc0cc519",
      x"38dd8465389657f884559362c0dca851924b9f513ba962939ac0118a9995f498",
      x"c57518a190785423828ef7cacc5c3cedebd483739a983b9e239f841acde952ee",
      x"373ac1ff526cc559deef357ba6e31152c378e5d4847155384b8791d0211de6b4",
      x"2237d9b37274d756e2e93cabe87510346685d195f2e7f4ccbf6b1fd74df46db4",
      x"2ea08682e8daed01e373b306ab2743d7020419ee2cd0d005d18d6fdbcda133dd",
      x"ac5ee17674bb1b9cb66ec22aa08380fb66908914415b99628a631fc318de3d29"
    ),
    (
      x"d4f9cddd478d9c400aa9294bd8faa569ecba472f9cb4c40e08224ebf38d59beb",
      x"44d571010eef8baccaa1bf0aea3b69b3c54d2aab7553adaf3d111c7db7a6e991",
      x"8bc836ffcb3c00d1abb8359a2b6280050217d704431f3ecdfc5cd1774f789b38",
      x"3eccd39ed85781307a4358d6c9731c420bc1e0003e7f7be50f5e7d81451599f8",
      x"7a2ccd44200e9fe4988fab3baa13abcdc4601727fe6e0c67fe055795a973e542",
      x"03d2e3a2631739ad642932c1b4d0030b7a335d332aa785f5b600dec7013f60ae",
      x"49c38ce15c69e74d38012b6a8d89e13993850b8494f50e4bb0fe4eb13683383e",
      x"d01dfba14952a91d2561d46d288134ca179232490ee40de214aebefaba020cc1",
      x"1f28f8170632bca7c3bc229bed6d3a710c308ebcfe1e9501c4244bdbb8387920",
      x"8f8728692cd959743dac8debb2d4bf66969423b0a7e158c4b85eac85a49d217f",
      x"90818faa2e6dc71750102d5e3de348200b56b8b1cbc70b13346b7a83c7adf089",
      x"5fd9a57dc3893d98006f54d56ead15460ca517970f80c7c99c40194d696f685d",
      x"90f17cd404b2d85d97c64ec9278714f4c0f23392773015a0db3ab56a093792a7",
      x"ee6188b511decc39202312efea369219e8c7e77db6f5f1cab230d2cc744e129d",
      x"20884b2603762069b42dd5a712b0bbd447c7503a00fe736aca5b8c08fe0cce9e",
      x"307279fe1247b41b29b0892248ef2a727a8c2d8bbcc6987d5889c9c5603a3a02",
      x"6a3df7563d16b1c5b1decca39e81f787372283a03e79a770a88aaa3e58ac13f8",
      x"78df75efc66cb75295e10d7252335ada87236ffe403567d83b295ee2d221fb2f",
      x"a94306101d784817d1d97332aaa7150321112aa1cacd40733bd1b837a991388f",
      x"fad732690f9bb7710e70c6b52934eb116862e3b5ee49746a4171bb9941827634",
      x"ca18ca7e49956a5e736eab64ae433f9cd7141f1aa05bb9d07c216a9fcf3e242e",
      x"5ae49c145472c0951728a2cdcd75f449ae2a22ed6bf96b4adde34a8935db6b44",
      x"0047fdb23dc368b2ddd49b92cb85202100ff0f7e5575ebeab9aae494ca7731ec",
      x"42642c5bfee5971e29ffb38cca2ce93a1df880f7601fef34be683d77cce76f13",
      x"f3cdc51c6e45bc93cf6bf0c84aa5b83e57017daa8a22369d8f18d45265694adc",
      x"88625208063c1ed6bfd8edfcf0ce636aaebb75837052e040d71cb21f562af1c4",
      x"53176f118ae427a3a0bad1bec8fbf989cb845ce6eb54f78a4a1dd25b4135d3e9",
      x"b1bd6177088d65d823fd9e2f7245f18a0223a0aa370c4b4a37ac89c55d5e06e6",
      x"cb3c85f59af8eae66c5eb23933a73ffadc12db38a62731e53111a419efb993a7",
      x"035e89c237fc5b432b54fa6ddadd148b13403f461d3da8ab1389830c00d09332"
    ),
    (
      x"6014ee15ecc62201bd6c1cf9531cfb4aab7551d5d265ddc6146d4239b763064f",
      x"490fd2cf1e167ac89f82a08f2a96bd15efaf17a6ba7e13b192cc9e03bba21909",
      x"3e21a91129566c1de3b40ad96b9fb9945e3641a5e79d9e087352670d56360aaa",
      x"2b847c2bc0fded99f53f82d06783936ce16a549ba9a400a577bd23c1b20de24e",
      x"815d75fc80bdf7012f18c15e5abda251969628b054ea99499b06600737ff472e",
      x"db3209037f342c0a2bc1ef75c5468b8f09a7249de1c1b5ec373c9ea27e3a092b",
      x"9ee56dfcc4d510c6691744a2a6b4f2e181994930ef395297b930801fd2ab28d9",
      x"d546e0427a10e2d2455e5610c8c42874a82280b769362e517e7265824a801310",
      x"9070f9c1eec4da75f4c578c7d168f1898743cc241e0ef04b6be98a0ef547a4eb",
      x"9a5053202878e1ceedd9631338481a6711e8bd1268967249bcf26b06040d5443",
      x"c918d6fd0994b4eec033aa9d5a2b86fb00f4347861f3bc2c92457b2dfee0586c",
      x"f4e2110eb95b5032a49580dcf0e005465dbb8684cdd76a14bce41f007d6a5bf7",
      x"99de6916504c9f3a581470b41855a531b29c7a5b4bfee9767f83d91c58c2e1ae",
      x"c28be3e0446c535e74ae1da45ec7ef6a9520f5787ebf49a8d7d7f7fbde058c34",
      x"9ae110c9e8c407094db8088738a6ae47b53b08b05bc276719f56271622c621f7",
      x"9f64ce0b35fa565efa28ec4897dfa65d7c3370262d6ff4422c77f8c8dc5000a7",
      x"956beff3d1c3d07220fe3b6b73a79ed00e4a8bd597be0122b63fa1cd50dd21e3",
      x"74bb1f3fb052767e672934b6d27e5f8c88ddff3ff5d1feb2486d425eee6f82b4",
      x"4a1192bd2269f916beb47ff3dcc701f3e48069be6d0282ea1902ffbce418f089",
      x"0ca529452a86ce4fb9cc82b4b3a9d4e9a23d395f01ffc6e596bcf1b648a339e4",
      x"7f84e0079f9cdfe083e0eb9d920bc1b09ad0ed76a344ea2c63b904ea274d2956",
      x"63567c209e939141b0a3c1e870fcb21eb6f49301ed26daead206bacdcd370f9e",
      x"8412d180a03076dd3b97ecd85f8154d0135be1f956bae98fa7d8896bf6291913",
      x"112757d5f5b1ab08529fb99405d229ca7dcdd093d5a04b0a2bb9f7f99e76bc18",
      x"d064ff6dcaede8b1fda96bba2fe6fe9f1717f9dc413f53b59d45f2428280126f",
      x"c427a83cb8c82b7356a059ff5658a86895d3effa7f8fcb93d916c4e99871f693",
      x"40afd9ad40a5d473145394bc938db405c7904de658655d36d0ef6e9268035584",
      x"1cddc0fe30e9a59a0155279fde6450109056f514ad21751ebc998a43ddac6d49",
      x"5c71f89849b60b8fc2421b93f861d21b225be060a90e7cf14f92836f78077cce",
      x"5e96c08055f417c17559bb404eb1825e25e1c7268f1ddf99452d44b5a5b8d43f"
    ),
    (
      x"1339e02df46f7055370653aacc4591c7a7496d916ab3906b8c818eb1136a4902",
      x"a4377fd9e92fb5df2459ce9a180bc990d3c2fff5c29447eda9cd6fbd1fbef56d",
      x"350736d5f1eb0c6787f894862ea7dc9ce834bb214af509b93f283a1f89e20e44",
      x"526f084a736493fd265815a8b6e2a2d844e7311add6e142ec48604d4ee0f98c8",
      x"5d802a04be976677a8b84d15505e747e71f18339bba4b72da7f34e168644309d",
      x"2b91626d51218f77feb3c5f164bb64c4b87f6c9c40bf2aba2a92cd9233ada541",
      x"ca0a5b7a326f7da742aa87429cc494831169e4c19126d72eaf83eba360dcf0d4",
      x"01bfd3f6aced3206db6f2cc23124e0bf49bc0f8e3e8c35c0277022364782a052",
      x"9923b53699518232967ade5b83eacd7b1fa31157556a8c4e2efed56212015b5b",
      x"8001d5236c2ad7d2b76acc9bbe16b2bb1dbed7268679fe182bc67803a218a73b",
      x"d1bbaa2d396ff13a9959de3dba7b5e4402f18c95790ddb4794514c5199ab144f",
      x"1879c739eb6c16cf7623c552fd0299a9de0e755f16d6b5dc1728c2cf25e0e82f",
      x"e840ec721f7021a50652a0eb44af928fcd63356299c6abd4665ff43c3bac8d90",
      x"eb3b9e969c1de3caf89d4f45918c8662aef8bb8fb8391ca5a877ab589ee4020b",
      x"48822c4e7384e6e6971a3e6c30dde9760e19f3e83bb2191db0ded9b89a934788",
      x"5db905e7daa209dd1936e18c77780628a971379c2c485174977dd67a60de3054",
      x"4a35dacb49bb0ed9dbc4cd1d9c5fe62c3534af85ec0709894e7cbeb056165d52",
      x"94d8e5d222470a9e3f1681ade18d2ffec9264247f6f9ae955704d62ca47e4b76",
      x"eda7735286a489607bb811d2c682a187fe5c6661f218e512cf0e60c7bb768241",
      x"63481776b95709df2c0f334f12e63e2ac1ee357ecfb05c23bd539e8509b0ce6d",
      x"8f506240a07ad4e724c50b5ab9cc421bdb6cb03e16415bc3a497156a4335b9b4",
      x"f864384506d6161831cda6b928d4524905b798fbc9351068de5cc84d0fa98145",
      x"7cd16bfb417590b8fd151df9c9fbd9f89c65679cc97a1a27bf1269ffac041bb9",
      x"1587de0f4f9f491b543a98f2eeda9b94945367c8a6ca419618ab8edb56becf84",
      x"6a738fac9385dcadded0f22c5f27cd8ba19c608c519cae50a11c08a9149d3fa6",
      x"88e4a681ac206d1b360703dea0eb9e45a946bae7d844bd52400f818130e05728",
      x"615e5afe959cc6d114ddbe83051d3a37f285a9033e5f60e0750e1ffcb75854a6",
      x"83d2cb22b0549efa9b499009a2067ee03582c4950ce2b4cdcdef3117aeafad63",
      x"42ee2c13d948fb7d0769dcfc5a57f085b532c7d6f2283ac915fcacd9463033ef",
      x"d4e8ba620143948ea6c51a06a2faab52dc9775d8a78cacf484f4024c3f4cdfe8"
    ),
    (
      x"498a2ec9f42b695686ea9e680889679ee5d80af570499ba8610f12e99e1b521c",
      x"8e3bed05a4c5955dc18e9244033d16cf8584d0c006fd326d40902bb11d91e889",
      x"9b75cd949ced806e8abc48b75a92bd2dea973334d32f7ae301b8fcd6bcc6f223",
      x"006b8e8935fee49548953cbfa52b61841e05ca2001923411fa371dd0441dc73d",
      x"0cdcc53de68b01d310fa688fa604ae6ade5be28604a583d4d8597e10244ace33",
      x"318708392dac9e3edba8791091ad12b609a3a44adfcca3bcebd8fd38625b43f1",
      x"c47296ad7ea2415eaaac7ea83ac3814a32f69076ad8b0e07445e023f2b3c3fbe",
      x"3de7ea043b86b534ab29390131d28fb73c7f0c837ab43e1e9d3941513e9e1eb4",
      x"512e3b470bd1e331fbdfa5a56eaae547206d4fcd557b329e75ee3a66143c7faf",
      x"6397ee4fe889c3d91c91b25b5d192ee2342478868a89eea98034066d7c87c683",
      x"e67d85849efa6c4ebebe0d05fa354b1b117b5ef3a5ad9880579332055bd33ec7",
      x"5c7485cb85983a199358018263ec3e5781baf1f95c113d08109f2933f3e26768",
      x"c45a9d29f17bc314f2356e38d894b92299b6055f429d6c53c198e323e1dca201",
      x"37dccd4ddf1990355534734270cd476bd6ca19d3e2d7e41781e825ee02565e66",
      x"c4f72a45fd545c48e429c88895dd92889d7d57bba29ce3fce2ef0a124a6020b9",
      x"eedd152d8db959b65d81f5cd3952abc239f83abe489226c91641d57109af297e",
      x"dbec477ae4ec9350ed37731584811b9da7aa933a30ee5e8a18df604cf3b180d1",
      x"bab7898b1307cf218d877f963782deeec4fc2d9d52a483f8335f45b5db2dc909",
      x"cdf45087ed00b31b14116b11edab59dd4b30b13299722fefb9fb6dea92c3c7eb",
      x"37c9b278392f0abe9aa9c8c8837ff5a8217c2d79d8d697c4d9dc170c81e7eaf0",
      x"77e3b8abfa90cfe61ac648e8c53bb222d2872dcf507b8efb58a8a7770c7d99ea",
      x"3c9bede8f96a1b2b4f9a46caab2859ebd270c5a816e6dd6312c40016d5cb9ad9",
      x"3ef09df260d7742d737d8de87daa852d14dda2840c0828c838269df7b13593ed",
      x"62a046c4fe6ed58721b379f5c31ac4bbf79253628c32aae4fc5f5f674964276f",
      x"a84ca07f515f802cabecbbfc8cebb1b2b234ed448ba424dcc81d22fa4ddc1e27",
      x"f324ac75d1c251c260da0b81eeea2a1dc9cf11d96a8cec91120caddc96999765",
      x"fa710635b77af156c9cca2bb12822c16b37f616c0bb2b097baca54acf8e982b7",
      x"5f0ea16b84be5dd09b43b447c531812a2bea7e6e4c93d6b4c1741817882e6ddf",
      x"d4f0e82e9e9f52c393a75898905e3544b1e1cd4476fadbaf02d038c105ef8d25",
      x"7df3c9fb9e70c137f103816e5538c319e973a6cf7b0d73fa9252cc27d995457d"
    ),
    (
      x"22c05106ae333c05e21aa2f89e145163dd30de5530b851ba6b36aefc321e64a0",
      x"fc0a6aac34545f1fc203bf893891ceed9e603bd47b2ecfb7bc6570b831f76d5d",
      x"a7658155cbdb877d6e2006bf46e1f1d8ba32137a4ae1d6087bcea07ca4d88314",
      x"833e05b0a915cd0094b880d6944b5be9ca18f6c3d70b391bc263fdd4807f1986",
      x"aba406e4225f45cf0d8b3107cf2a0a227cd26d1efed9456a5e5db6f7a52e6627",
      x"a36ecca344d71e478d6d254cc38f2640beec5a2a8b3d7482dc63bc9efef73aaa",
      x"66022899a3162f377ac78006af98800fb0a88e247450ced136fce6cbcada7e6d",
      x"cf6887da36c1c2457062255e32919f73b32e85fbd3c66ca777692be96f19a97a",
      x"b8e4ae606e8ab326d55b45e157a20f216b59935592d2386d6db02ebf60a3d19a",
      x"72ded81e39dbfb2e352a5716311d6b50561e842c118a8854a093f1dd620c9842",
      x"db2666360695b76fe31cb5c3258e3a307cc38cad584d72995f74dcd79b8539c3",
      x"1651e92093e8b302c82450673e12e89bf87b4d27ca1cb0c7a65c9a84ec11cac1",
      x"3adaa83ad1876ab7ff8d5002f947e2152b82017b0295ece86797192ab6799349",
      x"551120fa151c37c903ef7a467cbcdc5f6339a621ff9e56d1af85f805ecd40a4c",
      x"941a657d7f587043cd7fa99d3eb2c686ff52d0235050dfd6ceb1022e840de8ba",
      x"ed79a65992e1e0c1f75f5837db2e5ce4b0c56dce16c2bb93a80f311c677ac342",
      x"f987b273851e331778236242d0b0ef363d0bec0b75eaf3b2fc41b6ae74c85524",
      x"9ef09ec2d55ec4fac65bec26f1ac0c2bf70200f7aaf5904544f9ade59eb3c432",
      x"fe0b3ad954e163c0a66e3d52622aab252e714f0040ae45e9143fdc7b320b3d90",
      x"6a552c7350605abb028bcaf48c8fa1a5188fe417eeeef390b1520a1a59371dc9",
      x"686a43e7db558b3d62d5e5e6a4304e4db6068f76c0066bf75e3dc74d18eba2c1",
      x"7b966feed587efb41b6b58c86d5fd9f753ea2e176d125c4aa657d22af533f79a",
      x"f4f74f63d1cea75d5636ecec7823f44d532979a8dee33dacb1491c55f728e98a",
      x"8bd6fa8a9b1cb299e3b8136e79ab8a94782608d7b8f8f950fa0e490d6a94b7ee",
      x"87dc03fa4efde8aa4cbcf3f0121e79960d1a634be2462d3505c0bef88299613c",
      x"89207677fca69fd8fe3d3c8dda52d5f19c992c05644fa1fa96d4b076c6a04ff7",
      x"0af1fa9b142ac84105a842897235004b19e117079dc21f21b748ec36729a2b6d",
      x"21501910169b634a53058cbe534ebc8be744a77ae46cf1c2748ccb1a172bccea",
      x"328c2604943604f07fb4a0f1d5366f868bfbc99b1fcdc9f4bb57cbab95d60bf2",
      x"d82d9338a04361bc3d7c943bf266e11c9be3b70fb57e9d6f8083dfa28e4955b0"
    ),
    (
      x"2aa4d8fd425e6f2327025dc47703b167daf177aefa2851ff39158878668d76d9",
      x"e6770be40a0f0a11352556d8b685b5c545701418be670297b923287166e73ddf",
      x"563ee9bb701dee622db88a6f1e18363f539c7cc06ea53d0f5433283e4b962fa1",
      x"0b6e6d35afbb62af818e7d4bb4c426404adc99b7dc86444710659521d1d6f82a",
      x"aa0ef1dafa8d5479a8852fe801e075ddfc9df4f3e12cf5674ae419d2ddba3306",
      x"045ff3ba19cf8d09b862e8b9ce561f7773040879a105cf86f71364b58ab17e23",
      x"8485a82941f176599c64834a646c0fb853596223455e67d07eb631457e919bc6",
      x"dfecf5293dce71c0c8a63d989cfa3f70809c554516bd9a95cddf56f67bd76c82",
      x"ea86f53175a38dc827d4f178043b0bd4db30b4ce6dd2225e9a4c59a8ae90381e",
      x"974aee3299a1d1444260bd125b23f04cda4662faf90482406fec1fd15873a599",
      x"59cb0f08aa8a11a2c0c757c7737bc05bf1279c20731cd109ab7495fd0836e564",
      x"319171ef070a0664f8364d463ff5c0a10ef4d92996ee221ab72cb781e17d0c21",
      x"fb4e2a3011ea7be5e5ed6776f24219da6f0775d5acfd02de7052d1683c8b9a8a",
      x"2c2e8d2e15bb5f4b7031af3abb77b4e177a177da6cbb1d5932016af6dd243b2a",
      x"b34e31e16b00c4801f39d4627f853d2bd2b086c114b4022bcb4a04d8801dcbe4",
      x"4791abab59e7b5327c43ff852a0911cac33504b49832285ed75b50c3519bb825",
      x"c13081758ce9fbe0a11b7b0df3a5259e7347c431b8eb99aebaec63a5077b0a11",
      x"a48489c2c91e09dcfd5a1cff42161da10d0a854ae92e1f4668fb2e0078f36b2e",
      x"950640fd468f6e9985221fefa4f406dce5d4f8d0ca7737d2ea27d39d12625dc9",
      x"779f39437f26f1902fc3d0f2fa57dc2d3a4a73cff653c948637917f65812be25",
      x"5b8b37cbb3c71ab6f11be99f5f270886340ea74e43559065c77cb41502fc5feb",
      x"48c1c63e47de6c072b33d361d4520452076fcd4c52958446700e41d462273e18",
      x"28ec1789fde1497b91322ead92d725e66588e340cd3f2f8138d2f123be4ec20b",
      x"0591d056e638c060c58c9929510266311bc80fd1a73539200296a549aec56896",
      x"abc52fa7150c7e7fa905da5b806ac9f7bec43c8ca30ddd09298dbbff8dc031b5",
      x"0c986146eb6e0cef39a061816b4683e844a85d58da66b77f4301231848826157",
      x"c51aa573ee8cf4e2ef55a3a773f8902b9498b36bd9cbd88d81ca7698ab0ce99b",
      x"72595f95a92b0bbb3c0248048ac61a5aefd8642af6b4de37adcaf09330891cdb",
      x"ef8e39b2da080677877b0f255c5877c87d12719ffe73edcf7b50d2f10a7eca05",
      x"4a2008d667809bead4dde45d5d2a9f5e9fe3a44f117fc7069b3ae22b89bf2598"
    ),
    (
      x"24fda0c178f860d649d9be9ce51b27405fb62fc78721136353508b6c251c84c5",
      x"d6b30aad6595e30b6239ee75a6ee637b2671a2778067e348aff92d4317e2cadb",
      x"d4a93540e67200cf6bf416562f6314e0c877d7fab806aa71a6316fd3621c526d",
      x"869a8735e6b7b7975af455b76690fe09719b44413b1c08892b21c63f85c93ce9",
      x"021ab0e13c8b77f03d9a6b8160ef2f70f65792fe1c4fa0f3027c09baec347f5f",
      x"0ce1081ceeafea61996cbe71742e4af65b949ec9dde2e3f435687ec9a0c6ed77",
      x"cf336a75810da94c3c9bf9b954d22fea6a1e09f1de42c69d72a6cb3f5fc37d37",
      x"8e9bbbb721b70e64b57eacf382e52a16de8f6a21c81f0026eb99b6525804e14b",
      x"1c5286145f986ca68d2ee3563fc5199416dacb45739c4c6c6e390929a3812ff4",
      x"c2a0eeea48863a4a4a899b9a3340ff41aa6304b01a5e49acb9a5d83a4ec4b4a8",
      x"1f55954a51d92c5c55791c62a293d0ca89d2680c1fc251bcaaf5d5ceaeacf602",
      x"04ad9fe76e6cfd123531e8a91ee590812b99a295763136f8f14a77da8d6af4c5",
      x"33822350696af55862f81f59cc86ff9b98ff66d47bc9cecf5a8f35c720f90ebb",
      x"6b8099f3dce8ab0cfbd9fad93d075ba1bbac859753d19323e31c66e162865be2",
      x"1a6edb1efd9b42012f7047f0e9123683d8f268ff2ec42c4cbed736b9ce63b62e",
      x"f69633a5ee943840ef0c0ce15960a26b4170e8fc808ffca8b963adf1d5adf2ea",
      x"6b80ce6e37d37f8457481e81637d652f196e9dab9b3e6b9371ca5a6e4efa0f18",
      x"b22a3509051d3d32f7d03226a74f5c91a7ee91285a2a653abcb6e973a1354870",
      x"e9bb8585d2e2faf4c172a409bcdaf4eb1425a64d3f4afbd5137712f9c48875c7",
      x"7cca73ae3c4660404ae36f0c5fe4b49d6f860f45ddfaa460b87e42caa14bc30d",
      x"b4999ae06f2ab34606bbfbaa99809c1a36c0f5d50135288efac40c3f46957a99",
      x"0b6ac4be1f382df502d7a486de3bb1314245973cf71f6dd9d5e7edb1d0846918",
      x"ab98de55201eace670a669331ca00416c64b05b024e20569b152b0f6e6310af3",
      x"65d56cf9cb43ec6b06ae5da69660ce465f46c138800cbeaf85180e434483110b",
      x"3cf86f314b57e0de6044e3c6b1fb67b3c41e16ab1cd5dd9c94db18c7b34b40a8",
      x"24f17afc4d240ca7b7f87c77efd2590eecf18b0204638d31bf2b68b9752c4d32",
      x"58cec460ac75feadaae0f4892250af68311c75bc24219dbf4e86e69e908b3000",
      x"b62f3c878c849cd3202eb5c43af0ecdaa6f0695152082ff05402e0bda2432cd8",
      x"e87c433aa682f7b3bbaf3fb865096a67cf8b97e21d4f4329568bab1a4eb38523",
      x"1e8f929d6296a285b21ba8c8cdd1c8d991b456317f28e6f3f003128525a0015e"
    ),
    (
      x"7cc37787a4723e13e7a6825f3fae0ced3f6be1842c4df5000875edf8ab99f86f",
      x"64ef95ebe1e21db04bb756aeef166bd535c49f24899596fa6d7eaa4a3e7dbef5",
      x"8f81bfafb32af6af2feba2b7e14d10e20d8dd1b9118050220dd4fc987cdd7c01",
      x"6e10e69e8205e2691121a8ac3d9ff32be57d1e323de664ea4307a77d390ab76b",
      x"39d05a33bf4c46e12fd8983ab8d3b005e14da8472ea83f869902f58be9435b14",
      x"ae7419dd9872f001b3006d9d4440373101c217c2cd0060ae5035ba017909f5a3",
      x"4daf9d454af03f8d26b2e484d5c1db31df5142266a01db7a954506043e60d21d",
      x"a48dd379320172cd740ee3e9c6135da2d99005a41d42175c730ecaf8fb7090af",
      x"3071704d55565b9391190124a88fb195120b64acfbca93fe74a301bb6c8e86f4",
      x"3884728d5c5f3f976af19e2f9af07dadbd1e9b960dd6b391125a51f8828e753c",
      x"d84fc941c2e52412a2b8c1b313875b3d601850a121dfac94e5e2f2a0ef0e23f7",
      x"bad6c0e1a9fae8e49d65107fa91ef6f18c028b9aee8fc34eb6793c4733795597",
      x"99d2d3006d4a1a30681ff933d4de95bccc53125ba774d59f368e7d0fe8608f4f",
      x"182a4e85b002ec1dcd621644b707e51f9b4b4dd751789578c638274fc1dd07a4",
      x"bee657eb2a556c088286bd60999721b59939b459d871f412a43b6b4289ae281c",
      x"bc85d5d348c2f95e5172bdc4b632c0a3dc5a3b4d2df4b6098e3aec6e305bff07",
      x"e336d40c8ae018dd548000eebb98eecb1859626c615421c2149d84dd1a5be236",
      x"231d91ae29961e216f46cc43b3f3b52fd894dd795a206808e40823bbddf201dd",
      x"95c45755257693a0a3d8c0ba576e6a9e7c854cb9a722a22e68d6d97df74e63d5",
      x"cb4e79a43633cd475b12d894e3efe20a032c0de88e6532f59342ea6dec519633",
      x"e36bfae594727aedf33a19068f3a3b10f031fac48414c36c0812ae5272583e7e",
      x"023e4ebdc2218d8b7b6a5be91efc4db9c1b6e2329f0cccafe44c4f0d5fef85e9",
      x"a5c41a4e96aa72e5a6226556fcb377f60c23843af88ff72d3f09866183fedfb2",
      x"30f6943132fea55aee724da0a7678876f9fc5bed8c7821f773eb7e2945194389",
      x"625a642a6ba72f0a54e3f771e0c2348e9b30c93d4845e24269a883750234edd4",
      x"bdc8fbf0c715df3d5a3863aa9d8ae5b45499b5824cbe97238f2269d4fcac08b4",
      x"8fd7bb2f32cd624a5cb457a281790374e9a0ab9f1b92d9db7efd2e8fe9a4a66b",
      x"5f7b9b3c0859f4b71b60ac8aa388db0beaea312504331c77a953414affcd422b",
      x"49448a66befeedad5a0eb18bcec339b44ea66f6070bdcfd2849013255a1641da",
      x"44a694ea1d7929567a0d29d91cc7b8d617c190490ce8b57b589c915a505ad870"
    ),
    (
      x"792db055695b9ea1448a7aca82d44909308d316b746446d171bb031023699465",
      x"f7ba4ed58155870c4a560b26e6238bbaddadb7b86f88e3c07e06517c62cfec78",
      x"071657f854cf3c9a0d65c9a0bfc8b0aed354fd156b0e4600ce81bcb7467c3b64",
      x"920b92f5b7fd6875a32af9d6c03abeb073a26f119cb51a3597d34315b542408d",
      x"41b514d233ccf94f79a35b1582dae4656499419bd02f2f4f2a2339769a5325f1",
      x"fb5c68ee3f1e6270b4c2787a20a6484fda67254383e9444dcdeac931e6d1d568",
      x"fcf40b1c535c3f9a79eb072d66acc3e14f08198021d2128dcdad86257e77073f",
      x"07f12b2efa62fe62f47d85fbea245383fbc44d7ee9e0a76489cc9c29d5241f65",
      x"36b55f87adfdc15622771edc08f91e9052b49ee5a51026c7fc74c19fd249b6f2",
      x"3d47560c0ec037771cbad299ddea3d44ca452e173b5c623f2b1604faa4da2010",
      x"ff2e882b3de110b502974d3bc3f6046e01fc26e848f1841acba31f555c6760ab",
      x"b1bbb790a89df02ab0488154822d743bf51e0324540bfadd01387efac0775bc5",
      x"d9382f0d820afca512523ed4870ebcc0193e7a78569bef3dad1878d9f19e7f52",
      x"1982e7b9fe1740b6d199a12fe33775f1781491bab6e95cea5f6106f5369cd0b9",
      x"b6ff4351c290f85a1185e0787f7a8028e98934baf2a079bfc263e0f3940f2e1d",
      x"abdd7430c49667ed1fc9e5f2c5e4b4bcb0287d6fd4327820f37c15262317b7a3",
      x"d6f996c15b5875a1b43bacbff6660b6150e7d84e1ff6bef47fdb72c855b90690",
      x"2dd11d7d6439f41a3b786e75558cde5a2904b299afa0a9dfd748e95b206abfd1",
      x"f6da37ef61cf290b6d50bd9dc9abd1c52e15f0d38f0a52b6b9b2710353bff961",
      x"47a58d16c8fadfff1d731cea9dca0b0176b89469d1595076ba4f711f4950833f",
      x"c6fcb7f40ccc29563e7e54f5cb5b9b5b15d830309d41b57b03dff7549370ae62",
      x"f188c203e300953623176f85a88c507c4eef28969250ec0c3d22f951fb2149ac",
      x"ee177883964133a7e39dccff2af331cce4e7cea570f6bf94c04624606254d2ac",
      x"890615ff124617089d6fec34a767a155b59331adc0f4cc7b5885dc8354d0f6ff",
      x"72e6f9df3d6d0ca992524cde60e78f2c07e6fdae7a7871cd3c28588565c60808",
      x"6f313b4b3ec0a4c0f5230588588071cc4fb8c67258d515d617d1665885be48bc",
      x"3238880aa661dcf557d591ca5aa631905a14b2689a21aa8363f99940657e49cd",
      x"715d2724723fc39893ccef354696da5af05f736d4ee40fb926b060aa4ea766cd",
      x"2d16b900fb641386a102a5c4f33de42decb3fd9ddc8e1278627c88831690e660",
      x"38bf76b0b0c73c85465410f41e986020fb31ea32b0bfeb4d5184803e7107a4a2"
    ),
    (
      x"bbd12ca1578c52583fdb39218e134051f6e55a940d8c58b5a21665d85288e977",
      x"97b45e178dd2ddeb2a6ee980f15ff405489fea6c1616b3e076c9f342cb5956da",
      x"144349704882ec218b75ae408314720d2578497da38b0a753535e609b0b12e33",
      x"6f6f106586cfa42108999e8d462730379ea72b83a86366916d162ae0877aaa2d",
      x"0b4a9f63e6051ef68cb22c82e4e7be132c62123d24a8c272f1beb633ec9d767a",
      x"c3363a4f3d66dac18fca9535a12fef2afa651211e53b170b99590f521522fc71",
      x"d39d1ec42cd35b6f2a088c184c419c34fd07fc564494e36fa95dc0ea8e95997e",
      x"3a29e91c3b5f78d20ee0472d595a3e68c38ee5909bd6ac5c9b193b9f612fb14a",
      x"3291b68c8d0c1aaf658b826643fc6fc5d755231953a43697d225c31716cc8a5f",
      x"677a1bb2bf68f02f3c5f0d055209041abc90475e2d0f473ed0b648c9b882f5fd",
      x"1df74112320a220f505e66880c3518b6a2edd7988cde854620fc164b4f5e694f",
      x"442400d50ee88ecb7af90a59a1d2c153bd564c03754a472033771d34594fd162",
      x"e4bff68096f0e1fa7595858beb6732ff4ec21e97d826f4822d9d2a86a73f17a7",
      x"2152fe58fb012f7cf1c7b30fdc5b34d00665ede875721edfb0bf026927792127",
      x"b34bae62bca3c02503c52127ae30d853fce78a773040ecdf58a21d71f47933a6",
      x"d8cf8e56aa6baa9095011d06ab2232caef59251f6a93a55d53eee495f17ca474",
      x"2e05521281175e1be990a804f5d3e16c59d2b1171da28ce0691051fd0614d314",
      x"1c127ce7360a02762077c8d3b3c4fcaea73475341c5ce6bdc649b35cd00ae692",
      x"7a6db14a1f7e69da68b9b430e4ff21176c33cf0ef4e67a93f48a3d8f5caf4c23",
      x"95425fe609ea8bd50c882bb7c84c4d7ccebefb3a7caac2eb114df9c10cd00427",
      x"dc82e2d18777d1874d594cc3f0197cbb2562375002d0850f5b10eb047248b581",
      x"c76a997d256cdb8d2ab2fdb4e4afe4a415ab91adeb3b5518d0ff34aa531b73ad",
      x"5877ae28f0bb6802797ce8e1aeed09565f79dbb4500bfc0d2dacb63a1fdaafd0",
      x"3544bc0f773d5e4c4af9f8da835034228362840e44119c84f0dfd42b0bd55527",
      x"daadec46c27816e3623654905701b50fac5376cdb39c1c098e9f31106c461e3d",
      x"052212e4e0d8052a17ec2b1168cc60e4ded10d921fdbd7f60bbcbd397382d0f5",
      x"6ed50ad8d4722b3192078f2a1dcdcecbb86c235c70d7645c99b0c7f2da10116d",
      x"7e0ce356d434bd53cb2084954740b6ccccff72502fe0b8fcb531816ea5bf71ed",
      x"df2b2bf0326433d97a281966bd85be7041875a56b3c4a19b1bde8e0a198672cb",
      x"75604a97bd9da82661f479ca54f527bc00c222aa93a4c74907e3ded4dd6551e0"
    ),
    (
      x"4089767e649325891a1f1b212a11f7ce856dd34930bb858610046b14a66a0232",
      x"077760eb83da99341fa641346c5b1807e614e3e902491f972e97816f6bada765",
      x"95630b0ea49574c353d852d7067659357d0539eb9b5fe062b0ed0c92ac67684d",
      x"d16a5fc264f150c766e7b931a4a03c130d0f74b487221928ee8f953f224b2eb8",
      x"02a2fc5b8968a36cd85ce0aa2663238266c3e87b14b37ed9cd257113db536b3b",
      x"bf8cfa3ef1044ef53407cb69d7bc67ecb47fe6f5d6242411362c4149b1977baa",
      x"190a23980da5b93ef6ccff96733e1f8d3aafbe57e0017d883823e093517c3319",
      x"306a959ae226d16d510710b48e4f88b6104a3a0c566bab990cc5c4ecfaae5ae6",
      x"4f7762baa031b47e05c3d4aec17f0f4bec753cc7f166ef99ec7dea4e5295a843",
      x"9271aa27c1ff1ab08700076f43a95aeba76a0ba282463188c5941a957c1db210",
      x"b4de95f5c4ba9f4426bf5015d190cdd66ef1fbaaa4c9f4ef4ca0e3735507f379",
      x"6f370c322510bb1be5cedc40c9ca2e694c2b614ac2de0e582a94ad9ca7dfda58",
      x"44e8dbfadd5f4a876edd59d3894d11362af92fca87939312be1b73838e25d984",
      x"8c83126e49aa29acadabcd52a0fe1e3850d1484db17977e57ab401b8c44956e9",
      x"7df2b93317213780afb2a95abc755892fd41d5c9d7c8b3b28b9d02bb9aeb699a",
      x"304530eeb7fa8310349acf2d18fb9aad9d637b73d8e8860e3e9dcb7a1ead99e4",
      x"2a8d70f2d4fa9fa9fe27304424a4071f9a24d51ea267f32f5bce206e0e280a8e",
      x"6eabc44e65986913193c7ba591f82dbeadd5d65c3f85c7904378a3b53fb1d546",
      x"87b15d7fe02d107aa7a2aa529b88e66108fcb6fe1f9b9e89b933bec39aa2d61b",
      x"41eb46c01f7f41c8e5e3b4a3af9c1e3172b5595de1485da9697965bda088bf81",
      x"ddb3c15d7d743bc69a8f2027f04ee5f057e0bb1b973a5d278d7e7f4be051397d",
      x"9bff76e1eb2abc9495cee87acdd91e3eb02e6cae615effe0c6e833057254b572",
      x"1bd2e3d193e7508037af6d1219b94eb776b0fa3108ed1a19cb6a80adb2f2a4a3",
      x"4b03c62b72f0461d24975687932aac0efa884863da0bd28f23998215d0cede6f",
      x"5714edc661ea8e60c470eb156cf24863a70f2ce9a44f30f8b66f60f4a10757dd",
      x"015a841bf4bf2a6543fad9575a5821b20ca2590f5b366471952ffe8eee80044c",
      x"1189253c3630ecd97bd763b919321fcd86f6f8c3d27813e7a00480dc0da62b76",
      x"28777cff57f36125fb5af8e54328bd1475e30452a407aa9c4cdb68577d1f1483",
      x"081ce90cd1d2f1317528c59afbcef8bb157e81b43bbe17d4a4edf71243b269a1",
      x"0e5351ff04dd8a079666c099f4467449d61cea77b65e9c5a850fbc6719ad0c11"
    ),
    (
      x"97d997ff2915ad042c375ce47e074bf666f842c837a7df508d6ef576acf75192",
      x"9312d7988495263244a04315d8bd2b3ec1bb4cbbf30d9345a5bbef488a679839",
      x"9444bc46294ee91ed1140a0f1404a3d7a3a633215ccf0a06f9566429c613744f",
      x"2b54cb4a1fbb0d102ecd6be5e2382e0e1f8e9b277d87b5cbf1a3e5361ca1a952",
      x"41cba8d63149e8d7b3900ab514ebedd53e197d857991cb5d1750b16576400402",
      x"5132fef65a915ce0992e766895ca548843691dce309a4b398e2e689f8dc2f6fa",
      x"82c88cf090590873d41bfc442159fa445e8458fc909192804d397e0937b8bfb2",
      x"141a2d218e283c3cecb12542c8e11f01dedd687419f2a96f8a9cf67943d9c75f",
      x"e2ba80e7d83765c0c27891e5cc76d4966ae44a3f3409e2404f88a1839dd60147",
      x"0289bf85e3a46cc525e36e0923a95074c9e3b1bed6ad335ddcc8d7e7674ee714",
      x"a5711be12982a6ce18014d9bf75b0bc3e87d6aa23c5236af961b616a8b9a4663",
      x"6e11767c4eb5da2ff26935f8e9bbc913692163a3ffdfea7829b975545dc26a07",
      x"212f67c4be2fc59a55fb9c3411ac3e5259d10ac7862653c44cb6f9353e71466f",
      x"17fd0eea0bd8f362309d404ce9f13a80a21842a473b59d5d1eae7f3013bcb695",
      x"da4326721bb310f15ca3e0cde75af6f3c9a02598673cbea9c357bad2175b0169",
      x"ceb7a87c924aa8c9b10798abaec2cb5d490381a35487413f303d4a50a63ace2e",
      x"ba54d1a05c60a36abdcd3419f73aee45910f0565132b8e48edd792f0346dde63",
      x"56bc188644ef80475099d4af83a6b7ed2edb5e7d38e3bc0700dbb13eb46533a8",
      x"2f07106c4bc91324481083e492a8704ed4be1599ca968eab3dc5e87b74ae208e",
      x"cb47ed0db2f61161bb73f9531cf21d33e563a84ed054af93868b23ee89accac9",
      x"c5aaf81e040279cb30495c015d9b65254e187ad02776d9521871de9d25154c3d",
      x"12ecce31d116ea57c52711b369d14d88c721145d609a00f5545f8c858fd8d3fa",
      x"f56220025d38a38ce084a536b386653fd889eec25f9fda7452a6b229733b4641",
      x"b26d4deb7e162602ed1ffe1a417da22a8f17e73d663c08f1bfc82edbd65e4569",
      x"2af95be46e5368f61458074cb854129ea22d839efc5a134691231065978986e3",
      x"0fbe8605a0c5c447930592842532aae79716ee6d2d9dcb4e40acd0e257293a43",
      x"16a1d8d448484965c0ed9d037086488eeb8fcaf50799da6ad3906cd9e0d406db",
      x"9f0b30dd3f0a3f84cb8ce1c887842994c117acbe04c5584b1bc5759583008f31",
      x"1c269ca9c48c2a6720e3400aed686ae800ecbc7e770ce13df498e16895ceb2e2",
      x"dc4017ad4e42d304a965b38f4712778d44fa173a088cded19748ecc35c50e4d8"
    )
  );

  constant C0 : std_logic_vector(N - 1 downto 0) := (
      x"00000000809d4042d802e401d2796754c2f342290e3d7ea97c1b282f0dc8646b"
  );

  constant CONSTANTS : T_RS_MATRIX := (
      "110101001110001101010000111011",
      "100110101110111000000000100011",
      "011010001110110001110010001100",
      "011010100000101110000111110011",
      "100101010011010010101001100001",
      "000011011010011110001010111011",
      "001000000000100001001000001010",
      "100010111010100011111111010101",
      "111011010010000110100001100100",
      "100100011111001000100110111010",
      "011100000110010001000000000001",
      "100011111100010101111000000110",
      "100010101000001011000101001110",
      "100000100010100010000101100011",
      "101101011100111100010101000000",
      "000001000111000111001001101111",
      "011001100001010110011001000100",
      "011101011010010101000101011110",
      "100000000000001110111100100001",
      "111011101010000010000000000101",
      "110000001101001011001101100000",
      "100010000010001111111111111000",
      "010100000000010111100000101000",
      "000101000010100100000111111000",
      "110010101011011000110000001001",
      "011000111011011100111001101101",
      "101111011110100010001011001001",
      "111010011101100001100111010011",
      "011110100010000001111110010010",
      "010011011100010111100001101110",
      "000001110011110110001111010001",
      "100010011001110101001011001110",
      "101000101001101000010110010001",
      "000100101011000000010010101010",
      "011001111000101000101001011010",
      "101001010110101001110101000001",
      "101100100010110100111000011100",
      "101111100110011101010001011001"
  );

  constant ZMATRIX : T_ZMATRIX := (
    (
      x"8fcbf4e74311f40584e7352efb1803248c1959ca9247a9d07bf21d841e2cd20c",
      x"8a62542f624ea545ed178a5f19af246293f837828edd15621684036753a614de",
      x"1499c8a9bd7e8867545e3183072c06086dc5a32e1f793a4b8deef43b9189e3a4",
      x"aa8992983f7428e59cbd310a0e74d7a1575d31e568831b7dd245071e46124962",
      x"24d90d3935635cf5881c85e08a6cf0cbf3c09b4138874c754803b9b7ec877482",
      x"28d1753fb75ea8ce976ea4f3ab65b3fa274e79d08ca4e1f7c205ce02819684a0",
      x"78f6a113f21142b1d43d2351667fd79e5fa8428dff32b0f87f5011d5a7269cac",
      x"6e581f8e8eda4823db3769d57f50d2e2ccb8d00d36000c3d1abad444c3389874",
      x"f10a0519de2bb2d4ea1f711691c6e3df856f0238439084fa0000bb8193ab5be5",
      x"6c873e4ddbf416e41583987dc6fedf2802ee3b782071aa102025c4671ed40298",
      x"e57f12b6845345c3632713d0e2f09dee959e199641658a2ad94375610aa29b74",
      x"abbf0e5b49f2d4be436a101d748433ce5c5fdf8ebc7c327575d901dac50d4f53",
      x"16a7a5a8d3fc75b7d72932cf10dd6a63581ee6827979cc62620f5637714c2c6c",
      x"1522ff0b7320fda9b7c12e5103673a6cd378edd27cb69131ae157ee4826d8848",
      x"b6c714e154b4378237fb03e572dbe0b380c2cf36dea3ac37e3f62464a39c6028",
      x"3ab029c2158e156f7f63b0ed493352a3df6c35705ab4f3dd8c42d5b880a48ecb",
      x"7114b151813490b006de8c7b3f34dc7626bba7771c407a695db27bceb1bb11c3",
      x"2f0f2d86ef8b443855d630fab75ee77b7e10d1aa87d12e04313ba37e29c6190f",
      x"a8ce387c51a91bb2c4a0330607ba0e30d30486f502d5f8c52006b4f3084f57de",
      x"1f61e762f1896771926ce0dc0118c97fcd976d276642f7e8a7f3a83b15968e03",
      x"01c3929d693145db2da6a9bc6457a49af4113301084c595b1cd92d1d62195845",
      x"6e34dd4cd1a970db5c4950a3797702e220f65ec2b3e91429f6f78a263a89edd7",
      x"01618ce073aca3dd3c256801c67022f61b26e33405dff60b52b559f1b9857d9f",
      x"e1c69ec27020a9ccbc6bb736aa73de89b9ff59ae92809ac82781b68b070a6c19",
      x"f4b73573261a4ea79b66e85352966bb817fe252fecf594aa952b38b36dc454b4",
      x"c10ce703eac3720a23df1129b8e84383d2c79c3e69da0ae4888b78b655197710",
      x"910d34a9a1511f64ff53657787038481f79dfbe62f5929a5ad79d858b022ede4",
      x"69e052323f4380e3e92a65d0359d95df73c8bbaee4a74d8bc41523bf353ea55d",
      x"ed444206d485ff14508c8c8f1eed4f2671667e2b6c44541b38c415ba69605686",
      x"4b056980cd707ace501276029d7320d0ae452083a456d93dfd3d5044dec394a3"
    ),
    (
      x"5ee0e293c0374bbacbab516e2909d0aa26f5d84d600fc70ad11d34d5e740a866",
      x"9c88df8ccd87844d2d108e5d6f674f7b2c34956646840acead9229316db657fd",
      x"a3ba30f22908da1fbc1d9d472e307527e31eecd45532a81571f4dff69a9900d2",
      x"73e45f80fa530ef2b66f856d57648703f4482cfb23bb3ef7630c420a3cca5a81",
      x"12dd97a7373afd4bd83c12c0b2725825e1e29c955bfd7b4831f952800a468b8d",
      x"cdb26fa11bc9e5c209f8f8cb8be21bf39d30b11dd2d5332d9809c4a7957e0f63",
      x"b0623000894416486e84ecbc863bc2899fe17f050486c583832f4750077bd6d4",
      x"fc735af3f29db35558ed0ba8c4fc6af6a63b5bad5b8c20a2a1cac67a1723da9e",
      x"af8c54801aa99e30351a824969c76577ecf9b3d8c6c3fd7b0ebddaa3281819b4",
      x"c0d6e1824160b578d163bb40d841dfae995a2082281c064930b81c85bb514f3c",
      x"f85d802112426d9c1606cc7ca9653539ed79d6912f87f73c01428605f1472168",
      x"c8a935679cd1c41d0f645d0f076bf964e9e543186162571f4c02f1ff71e1a524",
      x"a30a2b19b4e93ea51e8afd4390b45a81fcd95bf3add10a4d9e9643299694a2f1",
      x"c8235f6ac4daa56cb2977d306ecdbd159c395ef54fcec79c21a08a0fde8c634d",
      x"130d4a88f597318fea7421ebcaade5675c9a8f0b61420291a16e3de841a6f6a9",
      x"596d921c996f5471c7800fd152deccb59a8d1ee3a035abded9aa9449404f513e",
      x"8e4ae6534c626df2143586df7ae378d13e0e91ab39ed157d7b94a10188d47a6e",
      x"03d20778d040e25d41e30e8aaaf1d3c72aa0fb8809043ad6f34b4a180c00f79a",
      x"086c69662f5f23a07d20f759a3fa8d69bd39b16be836f2ce41c767a2cc4f5328",
      x"abe65de0668135185eddbb6582d25ca8e1450e1491e7b292335fb787d4f85019",
      x"89efa611b025864656e7e1306d53e76a4bd98bfb5145c9f2057f60762b2e4f09",
      x"6ebbdd6ea7ef15437035c05d0938e93733f60936917925167fc0b52ba2956a1d",
      x"6fb2c5bf38051dc0bdd18e655b5f9adac91e5d6cb325a708cba7f1bb64735a27",
      x"06307093727a2741a1f9f1afa13e82dee0a0d6a2e0232f5a5cf8883bf6c99bc9",
      x"f53e08b78293d76299430f1cce57be22058f66247fd6049ba65b82f715429c50",
      x"0c396db4858301f2ffeb097a506612159760c2e1d86b488cb5e45453ec16b203",
      x"6aca640f28f28527d92cc7fc805049c688c42a877d6a77b8885af42bde49939b",
      x"2684ad107b43f9bbb95635a65514ad38f40f584e018140a6edddb4c67ae0f238",
      x"e55880b29ccc37f5ec840e796165a10b3e315874bdc84e5fa5ce7f4af31ac958",
      x"6ddcb8f37bb36e68dcf5a94f9f6f461cf1304c122963bafdb79dbf876cc4a0f7"
    ),
    (
      x"1815333a106a4c7b24a4d12fdf902c29a2c7b48b2db7cd9a0661dfaf0fe39749",
      x"035f429235feb9bf89eb6ae520de65bff6ac0e8117bd846b7d72d3bc40022b23",
      x"390281b5c8ebf90705aa8e81e8da62c55762dbc42c6720bfe69fb420d3ae665a",
      x"e22afb55095f1e507de38d3adc7070add5f902029823e9139d95f3ecb021b2c5",
      x"e1605446930f861edcc7eaa8d5a16d7b2dbfdb52cbc988597a120fe0bd2bc10f",
      x"8376a950aa5a723ae60663da8f23990fa57d22edbd641f084b47c7cedb26ee3b",
      x"20f4cbb7b3feab312ca7569b429045d55127b9fdd823e351abac0806c20d75b7",
      x"8bd192d547c5ede634f2aaaa3aad263de6dcb3f93feeafdaa33b032470d7a255",
      x"a2853c6433833f1f7fb2c3940928cc11660852473ba71ef23dace93785bb0b2d",
      x"ee4ea694fc68e931689b3b36683137feb41098e68bf8bcd1a7485a9fcce8da8a",
      x"d6eed5db14b0ed1cf5754bd195a8ffb476b3becbde9aa9c0b35d2282534d0053",
      x"59acdc0cc0d595d771419612a1a5c755a0ca844471c9314a1bcf377eb75571fa",
      x"eba55f5491fad407a36c394230c5f4a1f3731cab22a72a4bfc9cf163a6fa3d0d",
      x"d7dfaf3b09bc8f3126c5b97cc316611619533a1768baecec2e2154eea4a89781",
      x"10459758034fcca107df4e167fdf1f310f772eef343a14c35337ff3a85b076cb",
      x"c9256377b9b5dcf94051013a905e302b82e629d31ee93a6f104301129dd62cb4",
      x"9442fde04a48a522e5e95f257ca66921293f5e87ee8710731d0be1bb30b604ca",
      x"a797dc3121d62c39af65f532a2ffba7c0c8122e0d01c802db7088398da5ad2af",
      x"40aa4ccefe5a7a768450595c377f8b7b0c2416ff902067d4b9d1c16f19d6c40b",
      x"2317d2ba179bd8f05fb82e7725c42b7e0df64e186e5aa8d16809d874173fe507",
      x"14f72a5d8d4d804898acaa8a6c783477c973335e5b3ddc43447e686f8eeb1bc9",
      x"38aa769ed47c9f82ed595e336473a4df30e9814f95ebe5ef06b28fa681ae9630",
      x"be44f5fa8de7126942f1d2b947ed63f664226eaea78d6eaddb5096c930fa0fbc",
      x"5d0a069e5508807593d8138b90fc46b1646c33c0c8e42bc5f911d7969a90df60",
      x"14e95ac2ca4cf3f417cd674a921bb4cb5ca0fd3bb1c9f6c5368a839a5af98580",
      x"3b43b93a6ae307507de9b5203733e0b47dc2a78cf3df18106a241c067123e7ce",
      x"e25e0082e76deeed6c1d5cbc81fa172d02e1b7ccc9ca54c6b81eef893f4db568",
      x"6d054e6a1baeea835b837e47807ad88c65cb6e244f6ca08a8ed6329d40dd63d8",
      x"58d16dba0417f944eeaa88e5515d22065ea4ec4aeadadc1504100a0e360301fb",
      x"29baca6ce2c8f3e101fea116165d295fce315c2771926a5ca0792ac06f4c686f"
    ),
    (
      x"41fc3bcdb3eccc1804118c562e31d1649ccb0b89dc3ee292452beeb68380f83d",
      x"4d957aff9a62beaa570d2538137b18ff37faa391a95306dbc498c3bbfdbc3a67",
      x"508571dd279a697d599fdfbb729a95bd3a14ee700ff770b7f2b2d91aaa4c831b",
      x"2f08ebe419dafe8e8a0132ad960d2dfecc45dbd0fd59f7e8ac2178a92cdb448b",
      x"5533ae2a1e061da310f1245d0df08b4295f4439ac14e2ef9c78ed915979a14d9",
      x"545c633f4949380315367bb0df0da0d623c21ea0896f935043897f67ab61b909",
      x"e0528f27e0882d3a9a446a4c6cbcdc31f243687fe1d4d3a6cf31dfa21a6e62ae",
      x"e4f2091633bd6be44807df06589c96121f873409542abafa298ecedf6487ee14",
      x"a8eafd7ff05cc6745fc8121d471bacc5319b142a443f31a6f400a976720f5c4e",
      x"6205bb0fde61c25d2c252714007736dd228e7a8679dde0b7f4c4ef805a456b01",
      x"3504fa04d3b0ea53c8cb07e8d52d64cb60fc6784dbfa8168f80be9c403096665",
      x"5ddbf930d8c3ed7426047d68f8d913bbded7e623f70c673080c44627cc5c1d90",
      x"bf2551d25586a01921fa10f35d5fa4ac52ceec300133b9bfa26095dada4a02c7",
      x"08deca09964e990d84aa3bb0cd720fca2ea9c5a5e37c1be06f2fa2659a7935d8",
      x"8ff89e692ea3dcf0840bedf80eaed9e7488116ed92738f2b94d81ad5c4d9f68f",
      x"3b11716118a6ab4e77b87c021fef0a8616b89848ee1948f4f576fc629e72c1f1",
      x"3eee184aeb209e12c0e3cd8f63bf31d3e22215991070d896ed6547fa37ac6f5d",
      x"bac3422270f6db8c49437bdfba4e808586b6841d66162a61df51068f625070ab",
      x"c046cba020bbcc21fb1cb9acf68ad5503c73df89f343bb75bfa18e0e6f25e983",
      x"1fa995b749b7ab1b7c814ce92543c37ccac6447fd06bdb64df0659e8270d4deb",
      x"00fdd3355bed55b444122e0c1be78394dde1f99a4f5d87eebc081fce51ce3dfa",
      x"b1ba183741f13d44303104f7be9b9f4613859f863260ab7b941078c7943f360e",
      x"a0ac4e5ae3ee3c855c89596e7d42651cfc86a66d8b0351b60e276427da993130",
      x"7a2f049151fc5efba6b36cf8f2377a6a48d508303a9693a67b75e1d34a5754e1",
      x"b83ac3c45984a86b7936e8320b91f1d4a523dc08264e0ec71939e81e3883bba8",
      x"b1537bf6bf2b774f7fb692494584aad8fb7bb14177c4da311afaa0c8edc9e8e2",
      x"6c24a4ada9c7511db1b35ce093e313c09e61b90a5f61b2af1291285dbef5a181",
      x"76c25e9019a9439c5100f704a0d3a2bb689eeed21512a27edc2d50a7a215efdc",
      x"c302fbcad90aa63f4d920b11f7b83ce0653043aaf5702cbf3564570eb15070cb",
      x"7feeaf5f058d841d1798207c241a91ff1dc0597ec11ec8baa5cc79d34c194efb"
    ),
    (
      x"7086af8e21724d647252be55db1399e5a7a8bdf9fa8c9fc35ba75d668cd8a1e4",
      x"3592700595d69faa0b6d92cfd21044a3ed75b5a1361ed4a49c7045e41a48cc22",
      x"ed0685f6c5d8e56a41a93f9e36acf8a297e7947a4b193fb8d251c11d8aadb1c2",
      x"de47687dc4730dfcd232ef751687cb488b392dfe0861e11c64a22a35e6d24aa1",
      x"aaa41613f218ffafb023a2956adfa2bf618a4c9f7aee6d052fe19c2ac3ad6cae",
      x"a5f5c5d7039bc4ef9752862443915482d55ddc474df35c03b129c67844448614",
      x"5b1a1f794535c18c3a3d4b693031806dc3ffe05a98767eed94a763886f3e15e8",
      x"b62998dbc1ea47ff52979dde83b48b485ade6e116cbb4fa6e3fe573674c6b7a3",
      x"a755ce14b6373b0de4ccddd4db5cfe003f2164bfc16581412a1e69a65f47bc27",
      x"b3654bb45c73e4306f21a0eb7cc18b2f8d8385f8ebc7d1c721faed9b4b61a216",
      x"42f4f74e6532f2032dc7f8b66f23ffab7a1ce7b16d35ff5a7285e00c781bf8de",
      x"1de18f66652b332dc84e78688d83d9d9441e93550154f082883bf78519dfd5e4",
      x"a7f3f50d9f3c6a953ff492effa895af13774e6aad227255011fcaaea8e458ee5",
      x"ae3ad23c72494741798068d18d407280a0d457de2f01ee543d1faa26af27dc23",
      x"2efbbfed3f9e489506b588a42a05206c2bf0c9cf6c48347f51b80a3a0d5e4ee4",
      x"d7a4175241882b4cce016f7ea0b24413d322d846b78407c9121522a0cfb04f55",
      x"08edc75bccc6a1e3906bc360061d5cea91d9f7a32ffd0614873389dc0794711b",
      x"a37b50a700a9c744b9a66baf6d1ca4984611201d6485b08e1a2eb0ac237f0617",
      x"0bc4b6c2f80b073837a7c597e8c8a25a12479c37424ab20ee59cf28113e87590",
      x"4635faf67fe69a4ed7278389806112a131832a594fbcb2e4cf1a372e2d5b3788",
      x"b2bc420d2b136e66090b518378f956bb306a0f811b43c981528f2adb8d404647",
      x"a875794c01ad6eee8400219b81af89a4c5d8d6f8540739632ddf1f92be80f3a6",
      x"290680ca43f0a98ad7a5c0a6787bb40986bdebe47718308255fcedc2801568fc",
      x"19de7cf19323e44c51236e0cc245b3b9ea92f9b83bb86bf166cef1aa2c8e9bc9",
      x"b5d156a20225a626e1af847eade62fb6727edf005614da39d178f5a355e29003",
      x"0d4aad710ac0f3f25d106392fc88db8db0b9703af4dbc25216c47826cbabda5c",
      x"0f45c22e697616261b017f1ca14ce3d4d27bb33eacde3036359237cee5215b63",
      x"68d86c9a29f11f1fbe716f10ee055264977dcf3db60732deb8680e74de8e979f",
      x"e40e1fbc66d05d115415bd4666966861daff92fb4690fec9c9ccb50bf60d842d",
      x"5101e09a56da62fb68c02e64a326932aafb1aa006bc68ceb4fa3dfb35e51b98b"
    ),
    (
      x"7c2ff1ade2fb701c9cdac047c14e9514693e68967950ed7cb71e18a300a6cc8a",
      x"70f39395dac9b9a393ef833960b51aad67d716e8cbe03a4283afc39e79335a0d",
      x"aa025a9708e8cb8b098c8e6e6b6d93324ba62c565b7c7c798cbf70b9ba5d8b6a",
      x"8a7a0ddaa8d8206c0e13910daa4d67cf835ec2d28796098740c67419e3d011db",
      x"ad2cb1baaa9c6ad839f929552dbf190c399c1615d6f850d677f9e3a96596e0c7",
      x"6c24d372bc3d1e225bdf1d5c3dff371445000f25452831383289be4916ac3950",
      x"6058abf3709c1ae0ee32e62e84275dc021b81d0004bb0b7b6dcdf5110b2069e7",
      x"b77dc97a8841d4f3629335cca4ab7597bb7bce178cfca32883c513231074a625",
      x"c49e271d554d58c3241167888bf53dea029b9793b0982ca929b6d403dc8bca2e",
      x"e2f960565caa2af13fe9dd78a08e69bec541788c132c71d531a8158b09c175da",
      x"3a69cc3bbfb24baab098c01f7a58b5957660c8cb575d26196400f98c5824cb92",
      x"e4021a93b21464c96a0517811de9b436b69ab9df923b9de3a01b16f1801164c4",
      x"17279d7c36d57b4d18b6e48b51448cbab0097aa644214da69592186a743bf01a",
      x"f491b4c60a43320b32ea09e8badd30f9854a6950e094c34313b7baf5cd44b63a",
      x"198c7b5336a551837b98cec313bab212f789f6d48e1f6f8e75b1b3acaa505873",
      x"078f2649e03f4e2dfe807befc5a182c440104244919694df2ca38d866db52c41",
      x"c559ccf57b84254cc571d16b9632c2b70de18fe5c5d6f3aab2c0af2011c90a81",
      x"82b1417ec397362582e694932edd2ad0c4ae0958249fa3066dee941d7353085c",
      x"e06d6371f59ae16a7439405dac48779dae11d5e3974bbba761a6781e91144d1e",
      x"933af040251ddaf2e55348d99dde16308b64e1b726a289de2ffde2371a601a2b",
      x"572204eca6d64b2771404464b046797995268b8aaa6a7f040afd9132252d0342",
      x"8d1d3fec53b69d5113c9fcd9b488ad786953638546cc673cfaf36962a75b2c22",
      x"725848fb45405910d2716ece932f08c9827cd2073356b0f10cb6ed1b140ed186",
      x"a0a158d8512377982cb6801f11bee354301e6e5e45ce11c366a3f6794ede4e3a",
      x"db06a2e8a2b1c6a72ff799bb7147bc0ccef33c3f8ebb02aa7754f323a6c43098",
      x"c4ff2ec95b572776b9bc1d2818e306322f5dd36f0eaabe8b42b72ead6d68959c",
      x"ae191d0a6004ff332474cb569fef535b47ddf461fa1ea8913403d9186f09600b",
      x"22b7ac2d6f90f54ab4bd730a7821cef539aafefcff2ce9dfa2b7a3659b428261",
      x"ff91afe3fcae9d7b709723a57e65b899ef6d948d1077e08f5c29e4ca6cf507e0",
      x"0befcf90ecef229f16858e19c4225bd8c91f34d8f9bdc86fe9b78c33053c9d5d"
    ),
    (
      x"1abd7a9e7058781f9e3b832fb28bda30f5756923190134f276be5b619df0af0b",
      x"97c7976f170fc497a86fd466da1d3da5ec0db11cd9ef6a115f941af0d980bef4",
      x"035baa7a0d127bcd2898eb61d0e3dc113144b581ef3c1cac5bc74674cd27ce2a",
      x"0934b1e5699321f1d94152287b708259ceebbedd3b68824e87ba279377a8e3ec",
      x"6871ff68c16e62a764a13cbc9b7b8c295d95ea8b55522fd3b8e0fb69605643e4",
      x"4774e4bcad5b8f264193afb2de262a7e998d2b645177ad512a69213001475a2f",
      x"08b471437261cbe74ed26b807127018a1a9437acee5ee3c80cc256981ff2d502",
      x"d16ac2745d75929969bbd834d3badd1dea6c45dbe05f2d99ac2171fdd9a680cd",
      x"2cd01db47a8fdd598db3688d1d0650e3498fb4839318d790b04eaf37ef0514f4",
      x"9edf4fe4e21d5ceefc36fed927d2c6f3a8082e6d0615385a2961e6f08a1a3689",
      x"4d867405e40b41d99b1628d88ee89668ff20af6c01d6cb5b5edf622761f5e55b",
      x"1f4690faf307fc699773bb8ac0aaafba984019a45ab669fb4b91e9e9a2796579",
      x"793a6b1aac75b6cf7f144467692ecaa08969138ebf112e935563ce5bef810797",
      x"35cb6c73184950a593dfc4276e26b7446e756e922e6c56259e8886ce53ba2f11",
      x"c2f60a6472c2e7f5e9215ffb364596d9a9e8988e498a49e66e2a5780c794171f",
      x"4c027da05748a13704cf88386535db5287ed05f5c984a2d7209f8c19b0dbff24",
      x"eb64c0fb053da6e344d91e12ec5ca814958ee6bbb48bc7e561538511f4531cb7",
      x"9b902d2e56cb326bd52caef7b154434c74bca07e73ecbe2db1296b97d28551c2",
      x"fcfadc850bb7eae7febb2415f45b4850d708ed96ebfc0ee46ce5cdaf587734e2",
      x"2c287edcc189bfe3b602417aa4f58ebd4fd178667f5d9da0bfb684752319cf79",
      x"d589d67ee726c5bb794ac9b09ccebc792fa4f93bf9eeaa048ef348edcbb7742c",
      x"3facc0a6a8462952a31a4759d0cfe19fb8f633552f7616af5f368cf9a216c426",
      x"64cf81b9c4f09e35443162ba6df9365fe519bcf2ee9dc14136a3e4d412e6bec0",
      x"be092852d771108c5279f6234f42c28e5a66b25a19c50ccd62ab97a4c656e5cb",
      x"3c964faf87a4a6f30808e5298dd01582c3cc7368b36a4b82aa9aec13dc38749e",
      x"4acac94001d18040b095dddd826c789b0d249d879bb927b736e8ca426ac4f950",
      x"e3bbfe875f143058f793bf331bf952b256add6e56ddb57e1cf347c6ab34f8ff7",
      x"823b7f3bb906d873a081e5a85ab01347658fe4e04cc231c55db9ad9a33d7dab7",
      x"555a719f550e23f17f65d5e4955fae22278f7980d7b1554d9ca57b72cc5c853b",
      x"94baeb5298be44cdd64e3aa93c20339ba17c06d022fa9ca9cf77f4d1988b2567"
    ),
    (
      x"06f8fed1b37136612002ec0dea25d6a7c244326237e8cbc91572328720d68da2",
      x"1d24559f3618fbb6716635d057fdaddc1008de630758e9a7d0205e5f99792f6b",
      x"4a3bf24c190091db38eb606ad20d191c9a5e1b24b9cb286738df01d1f0af3704",
      x"972fb003f3923983a09a23c3667c1963c6aa199cffcde67053d51fd7d3fc0400",
      x"7096f6f8e11de5585a66de3f9a91f698bd8a1b17549314a10f900e481fbe98e4",
      x"a5ea55f0193fa4815304f2bdbd9a2cec5b12f3f7996cb12374fcbd69c63c1e96",
      x"4033aba7978d1f72dd87b246c551537caa35c52407cfae871ab90069181956a1",
      x"d93ebafe52b906b9f7bbb9930a0e1bd368623bccd965e5306a9ab47409442b46",
      x"a5bfde64ebabee59e338770067a54971b4950fc133e78978f42da79fde228fe7",
      x"6d1fc958bc0fdde932c4b9ad0c88179dac12bbb93055201395180f896c7471be",
      x"dc48689ae4eb07ee7096f8aa105b70593eecb4cdeb111d0432b1ebc744179e0e",
      x"36afb2a502689f26233997894c81bc4547a1d36d4e46098e0594030a351eda66",
      x"0c6b4979e9b2f5b26e9dc2da26722dc49c8c69e94a79e7e63a40c260ca39a97a",
      x"57ee31bd4817dd24b413134b5b796082d0fbadb3fad6721045dceee0e8104133",
      x"72cd34eff662b039b8f7f90a508cc2182e8ed15f86001f8b1fba707f6ba7c650",
      x"8a2e0d437ce1dfc1335b42d5f40298622f4b48f1eaefe6de8da4a0eeec420477",
      x"445c654200a382ae96ffaf763ab839614c96f73b6ca9e1cf1a233793260a694e",
      x"e4447b30d1982a16fa4a99403c9b06014e637e2b28e62fcc56b80630da61db00",
      x"74694ee10c52eacb566a277001c9e7a3a4de305c2a387e8afeb7362e5ce55644",
      x"32cd0d0a75983b1b6445095b4c3aee2b8a1c9108ff778c3568a9dd875d490862",
      x"1a20a7fbb05713b056201feaff4ecd895e9e6fa85824348c734101ae435eef1d",
      x"ff595f12286ce3f9c1e5173824c31167f9475862d69696d3eaf17bfcc69e522c",
      x"a822a81260d43d37da2ce44f65cccc1867c0888fc546005eb054c0ee8d3406b8",
      x"fafccbc9fbdea0e5de6c277e67279d61bebe4db94629865091eab35d12304476",
      x"25d35905fc9ef82aded4042bbbe0a17102b7f2fbd662860e666d7bfbbb760233",
      x"36bb9e4177486250fc5f75ca89ea578374c8508f74e23cb8b8d2c7d16a430a1a",
      x"39438a10785a29c5b4e6181e7c049fddd31a9a33bec5ee3e6f6f3ec9acf3ec05",
      x"1bd8f6c0b97ac7a4114028534c99f2b2b48f6d05803bd817882330b0a5516148",
      x"224fb9ca379ace70ecf4049360ea2b8a6eefa61b7bc2048676d014c1592dc3e6",
      x"c5fd4e3c4bd3667b30740ed57ddb3d05f6868c73c7aae9dbfb399c0cbf210778"
    ),
    (
      x"29467fdc4d3911bbb3a6887578d921bcb696e87d4b21ba6e106c8d81f70d16fb",
      x"9317a245634d39dba6eb56a191df30ee29a928ba5414929f6392aab3d485c45f",
      x"ea0ba1de442d186a9a276b11ffc0a95dd4a64385e672427e73a84665264ab8e7",
      x"9544a1588731e4f2db9276be447510ca40de3d1fa4c66710bb8c84eb3c4401a4",
      x"f8d666003ce609360b98f0cda8b029641c9f9010229347055408bc8dd6f17338",
      x"702aac3f4ee55d38827def7284488b4c95288c10d185bb175aeac4df05b11b45",
      x"9aead3f8759c6d75102686f68df041b660fb63c3819a6e939089ebdce8a61d68",
      x"ed234b7a16e74e88cfa3476ef620be028ff38445c39d162ec8afeca503098762",
      x"9998f98d28713a7c9f16df37560ab4cab24a7766f4937b1a0db4d6c61f2063a7",
      x"d8425dfcde8c45ffd2286a31d8818f252a19628f7b9d295b6c16d4fe6230d369",
      x"afa0800176c88f42aa63acd9903dc3fa0a2311ad5c11d1c7c629997fd51159dc",
      x"732cf7c4bc4228cd0d4f3c616250f13e4646d9931803f3e2212f5a30d2d26ecd",
      x"2b30ed8eab76f0cfa0b47872372911e47d934f0d2d759d8e9de4111d061ef584",
      x"307057ee770de8b95fc0270f693f0c7b5d062a264a29b33436831c81f81402db",
      x"aa216466f386bf946afaabe399b31baf9d93ed5c0897fed484fa2fb479bdbeb4",
      x"3341aa17178d6600e399f3819ff9da78084528b9418733b212a6ada4347fa8b5",
      x"262731f2d66395d966246d3423452a50bdb610f206376de0a278b3c5381c67c2",
      x"2d7a27138695d0fbae20b467eab2556b9e6560a3f486907fba7f3cb048703a57",
      x"cd370198494c4e6c665e8b6a5fa0cb1598f89be00d11cc58b3410d48e9574f7d",
      x"e40295169c5cd7088fc0c47b3b3a1d5e79ea3d8a0098ae4c3f52bdf443c8cb62",
      x"c9e4a609bd3a2d8b0c9f38f6f285cd8826ec18d9b945c84c84d4fd1f022c16b4",
      x"27c6550e1382d5345ecdac30ae2d4d33ea5ce6b8d741dc0ea21abe8f544ea458",
      x"44f8ef5787b981db10d507d7b0a846e45f0f126e226e3fe03cbf095eabaef648",
      x"7b990a27b6bfc7275e0be6da8c2f1daebf1900ae18a621c38d3e51b1bf0cbb1a",
      x"6ed2d6e831828ec6ae77fb0d64c12fa97f81028f7c9bfc944202b4045dd8d8bd",
      x"1a07d5534e1804b6cc1e7714d8810d5e938c2f1d1724dbbdb8ae17cde6aaa7c8",
      x"6e7aded0728de2711f2966fe3a6e9f053755a8fa62a5a48f03ef08a72ed31cc8",
      x"882838b4f19d28e6bccf9535d8eb131f461533e6ee22266e06d09dba8eb69399",
      x"b11df439a83843279a477da0cc545513b60a71552ba530d8e39ed5035f327d00",
      x"cb63864f4000e4c500fce5203b7d02c3141bb3ff25f0509768d9e001f76186b0"
    ),
    (
      x"ca12cf173a4fc93aaa3c70c2d16b414d5995fa07bd27ff06e534f61adf576da1",
      x"80c0a3ecf9ae4891ed6eb62539bcad346578ed4a247ecd227638eae58928af7f",
      x"283aa63fa8c9c24120a2592bb7ae30bade70dcc288546c4ffadbaeb7f5012c69",
      x"3d152005e22734aa42302913442c80051f9871593c6521275b98da62995676a7",
      x"f71bf7ef0cd3948edb41143d8c282f49000d8b0bfc62246476c9cd8b1c2483d0",
      x"82ae2b40807bb5e780ce0cb88c64d305355c89f44b4c1373d5a170c8c48a5f80",
      x"b291eed445d2df0974bf878750350eb1d75dfce7d1176086246a69657ce832de",
      x"5399cd08752ad9c55295e6708bd24720629330d298abfba63f2bbf5a7d865d5f",
      x"ddf090e40dba7fce63442a15b008a45b16068af17273a0d16cc07aba19675692",
      x"02ef3fe391e4449bfc9c9eb518ad22b7e152e8cd0ab990eec937effbd44258ba",
      x"17a7490c9246b98225f90505ca0e2632c186f980e6bb76800d0f9d5120729c41",
      x"597047bdb20e7eed4e248dbb719e76e11748397076655d6fc7a71348e827209c",
      x"d631865246fb73bf3e8960a3956b207a3aef1c6fd9db30942e9c5cc98744597c",
      x"923aa4f38a6e4f9872cd181d194e6b89f3367632ab2c8a3f31e0b6414ce94eb5",
      x"2f84484c92e70f6ce1235dbb91d4c4e7b5377f5ed4989199bf50df5a513245c9",
      x"b603f7472ff07b4cf04b7a8412f309dfe9cb0511a318e4324d7ef488fb659659",
      x"dcbd650aa35d6884dab34fcdd04e39d0af8d1746942fbe87f447e8ee7155584c",
      x"9ac79309305379e426f7348923c5164e142fb34aaae0476160428ce0ea626aa6",
      x"b40f78da5bbe061a5e01ae0893c4d7407b0ce0d18cad6714df0626cb776689f2",
      x"db719e5ca6809bbc17213294640b3a181111055e4853a421b866c8cd7371a51e",
      x"0a23cc30b613855a8400bad63ff953a264d079ed2f33fda0b8287328b49f1cc4",
      x"0164d39e49a9e8fa565da1f90324255ae8b146f4a61e4077133f7b1d1a2fb8f4",
      x"e43b3d6d968370ec4ee76830ac52200a0c837f287f848f17ef96f44f09aa5d85",
      x"31eed534810ad4795be24c0688768d9910c311004d44b0338d2564c2694669ec",
      x"45876b7d24aa088b2b65a0d8d48100842fb3d21759d00b6534d706b343c50f77",
      x"3f5afd90b47f9936b468d25685494f6efd6bf50ce49ccd7abdb60f53a6af5bf7",
      x"bdb9b4f91826d71383bc1eeaa2a9549fe696408c2a223d12af122ad4a0ae7e51",
      x"4c465e6a9126e5656cf5904bcab66ee6940519b50cdd1623d0b36e97a7988561",
      x"886481c8ecec4cf4f547f8a05bdfb9b2a3892f6b4fad4bda0e508fa7e50da714",
      x"5472575f3eb87670068fe6b07d868106872a84b2419112062c30f0337b5dfe62"
    ),
    (
      x"9994bc8f0e0d1e9f032867cb75d22fd53bacf71e06fb22e8dcb5b449e15ae60a",
      x"d1d1990379d788dec2d21add81aab2eb30aef0926e1a33b63cdf4f0989f3a8fb",
      x"cdc768246f02e3a909153103e957137e0e604986b91e13b370a47ca1e32be86a",
      x"96d9124bc755e06d885330f3f240622a2ffc6cdde6c0e489504ef8f064c2cda8",
      x"faee1db0b23b0b78799d78fb6b60141f8c738f070d56188bde057bc186df3cf2",
      x"2240ab224fea44ca762469925f2bbb85f9d79e34e1feefa5efbf54c682dc0ae4",
      x"96a7766d2b39a8630d64a022aeea7c29b7974bf509d4be17c8f4787feb88bd1c",
      x"9da3c936a3eaeed0ede61fde644330dccc8876f150607455d881749b2707cb09",
      x"7e9ec54d2e81f82d58d6c57ba3b6d8a65bdc1e4b57a0530ce7bf092bdbcd2be0",
      x"fb37b036211edc6d0076ec11713ca506d57a23777837e998130f8304b4ba5b42",
      x"c9356efb681e7aae14058758c89a2a1780be40638cfbf2dc685f7d9c49abc535",
      x"53665e493da2f37ac830273df1948354c49a121ad9104bef2369a97b9037bf66",
      x"a81d260931da9df61f67e235aeb6a8dea6efbf9d05c844ebeb510b7f90cb1d90",
      x"b717fdc6d90ae2705d96d53a9ab54015683e26eda83fb3128029c628897aa35a",
      x"8ebdf892114884d25276406bb0107b33ecceda5eac8ae770bacbe7d1007ee07b",
      x"51782921c8ddea82c6fff1c96373d408519953589d8f3f975556265331ccb865",
      x"acab58281fa130f5d8d3548dcd31e2163a3dc251793fe8cde50a689007e399b7",
      x"a44c05b08809fd2401dd0292dcbfb517354a1e3eb6874d4cd9377cfe9cad66a6",
      x"d6e14c79f343b86395b836d6a9cbcd16a254236333b5585a09c826203498c840",
      x"0523c3a1dc8c97bef3468308e80d521ca12a23ee3745bed4f86dfa652da4e052",
      x"42335e9977df68e3156fd55e7685fb1e7109a3f6570534b5dc094b778da30102",
      x"6f6566d34a7d400b690266d07ae2dfe62ccc2a9d242ded257086e6bf90fa6ec2",
      x"4ea3661b835c498958e7d0834f6312f8b69e0775d0bf309afc36acb875c664c6",
      x"061605cadc68d6da03755a7ce24e57b75be6fbb5c513c515f985817e36ff8ff4",
      x"b02f2e726257d7c61f4c127aed7d2d5f395887666b9105e2a65c8bc0a441eedb",
      x"6e4cc0268cc3e9c18202b21821b95e81c5b7b15e753077ac4fc493c7d08042b3",
      x"69ed0b1c786d6d05d395b570671d6c42ab3aabc9c88e9abee93872d9e3cbe053",
      x"8d68b8efa7895349900fa00a4a50b67d6aabc6cc4909da07d9d62530c9f68069",
      x"1654fdd1366abcdb480466d989208050e69177f7bb3f1e15f9025c8e49167393",
      x"db9bbb34eaea20be250ceb38de453820c3596ec85fdf6bb806eb4114619977bd"
    ),
    (
      x"9ab6c853d3a51c97711e21c77869301dcc1f51ac524c73b4579ba64fc7f8fe5a",
      x"9cf352426930d62bedca4d7d2725a43021d8ba978cea07a98051203d69667bbf",
      x"43ed95fba7b02bb22d12c2f935c06b72857b368b17a5e0e8adf724489f16e047",
      x"684942b397310981c86fe38302a1abc2cd0bf9cd033b917f12e0b0047210cbe5",
      x"50eb08f72bbcb4b3e06f2344fb69fc26fd074579264bb1f267b128083dcd108a",
      x"2799f3d1669d61012c5e493bbe0384cdab70c2235645332c47597faf1c2e6788",
      x"7bb0e2ee33252cbd5341ded50e82bfce6cd1fc56feab48a0cc1f66df35c56956",
      x"7af1552ddce7d7ef9f6c79d41734958b85cdf79f7cc234bb40de2cce2a2b8a90",
      x"465a7a7da4682fcd3315af46b71aa2bf7d4d0e4f607f74ece0f3446dd1682d11",
      x"4e804de996ca749dea0ba55a07976f59d4448ce3101f132d1d6e43802bd80aa5",
      x"17eabbbac9f4fabd21849e090327b54e7c6a599b5b31b72bec13949a07629913",
      x"b206c9e36594e6fe24cae76190f53022a4032ae153705ea89504bacdd058877f",
      x"dd34a77f7bca945e86701a3995d07fe2b243961c56df0250b8fa3995638eb282",
      x"ece3da86403f8ce393f97be4d04e56ea3b5772c4fb86e3aa54c9ffa517dd7195",
      x"65c56b201eee4e8722e2a44e058b5a39280cca75c301fae194af9cac755143af",
      x"cf2d87f4897da106f05b172a749c6a4c2573f820a4103a63d234f272dd1e5562",
      x"ae8f04e17d7b0313c5354e463b4156c11219f50a5f56b1f07570d4a715fddfc4",
      x"e9a35a1086485acdd511c1c5b8713b9b08d0b5a979e0800017ad78588fb90664",
      x"db22c43613ba6a122306fcebd0e114ba2c71c47ad313fbc550eb86e41bba99c6",
      x"658861a8aee6763b6561d263fccf5100384bc169327a594896d379dc0fd4f580",
      x"8fd0965f8b8eb22b5908b14cd05fd9f8c163a677afecbfb6104bc1505b345032",
      x"0802be334625f5de1ac1c69fc9ad7784c7a709286db6831c6e1838b956226b27",
      x"7bf7baccd187aa0bb0275fa40b86af507c15b4354f77b69dcc09101ec27ffdec",
      x"f2353383eb34010d2e49ae15f8c68e504ee89c126b631a5e42aa2dbfd29b7721",
      x"b695499bd1c034c4245cde1336ccc05d2e6a915ff19d279046d8280b8d37969a",
      x"8eec3e5cb78c5b858ca443b2772433ee87514a45a5aa45dfb1ffa60f9539ee05",
      x"74b7a82b111069acb1e9772fbc71fe7ab284674d72e055349961266d2427515c",
      x"d4a3c41cb99bb81e7f7845f2d3759b5a643afcfc2e5ab4dfac4d73792cea9b47",
      x"65976a3dbe1a1a1708457031da289500d49df6937f5f5b252ed056cb3e12244c",
      x"7dcf00848e233ad58fc295ce767974e63aa2a92870a895a94486f85ee23430db"
    ),
    (
      x"4db60607491d0d8a983e754d5f9c9536a001cbf44f15c1ec5549ab790777a7e8",
      x"1064bcd246de23d803e1c9eafa383d80238293544c1c5e25d1c8d90fedc98213",
      x"8c71c2af9342ccc985d644c825d950824b9e7a10e10d7df03cdd673536003316",
      x"db3d339baa005396f9e04282ed55395bc64c19f3646896b5679c979f009a4bdc",
      x"1de90feae674dc46b8730b22f63201d92ebba548cdc427c10c1d8924686d480a",
      x"48ec79e74692a8d6b553102813748c62e8e2073f6de192e2f522250323624259",
      x"e4629a3a4dd87a9be9077a41a70c57ca97c6ab06954120bb309ac2c94ce7b5ce",
      x"679c277eebddb248f04015539331c69071231471743eadb718cc352530699a8b",
      x"80745d4912f0317f3ca3e53a66dd895078cd42fb3909cd3e39a3999e843eb950",
      x"e84c0e3cc30e6a1619a5df99e023752cfc6625b873b8817444f85587ad3c51a4",
      x"b4c806b21b4a1abdd033a55942cc45fe64bad87ff5b710f752e1c82fcd7cf8aa",
      x"38767e328a29743e7582a6935970848856fb1dd53ec62cf00db1f6f157214bc2",
      x"e16ee500f121b3d1e641f5791c9f907e54b39b3a5b777a605638e012a84f7785",
      x"d79e1a4f16980347773fe7361898ce47d109a4246399be7cda12911dbce5af87",
      x"2eefa50b4f12bc946a3413de2079bbd85194fa310e4c9eacf3de18e4f0368a9d",
      x"cb388963c98de88c9aa65e92cb845e00f0917b026d0e273b0ff6c79d7f955fd7",
      x"9fb49a484b5ee88736722e0f23a63ed74259fcedbe70e2abdf3fc49c2110b68b",
      x"35d74dc34a7c90fa2b65b0392a22131f51a278ef7fc4f0c93bf25c251411fe8e",
      x"8705b1040b9755f8b92c49cd3d372fad3ca32bb2ae2fdd761a59b48ac930a5a3",
      x"3a4fd7091dfff70e5c2d3c434eb756100b1b585ce402b73f4874dc830fafe2a5",
      x"58e828d2ea77e43c043dcd1fc79c437b000a03fa15dbbc84b6b0f7ff7f1f22db",
      x"43ec12503fce66248377a6dfe8c83683aca453867fbe0c00c1a6f45d32b91d51",
      x"f86671dd475d8a0e80fd51b15925c3e18c8ec95cf9fe69b9a7558d94563be0e5",
      x"0c42c7fefca0733c557022caf901602a94bd6119317fc14524d59c72ff4b5dc5",
      x"55b0fe7563b672618a0e4f4c1ab909396b813c7c5c69e97353fc5710752b0497",
      x"08d0f1dd69eaf34ffbb4f5a64265dd459ad8ef699748c97a4884af2603ef50f9",
      x"9629feece9db3f4c16ea7d1a6fd46b7aa28a5547087cd8955afce388bbee16ae",
      x"f1b8f773ba04d8b2d055f0e7bd4f38845b66334621fa99335199c43077c28c90",
      x"e01bb93b949f1cfd304ab9bbe5c77dc3555369d8def143f17a77a75b8dfdb625",
      x"aa56706df8155df6f10606158dd5d1afd3cce10159c336cf7f0a0e5e57252f73"
    ),
    (
      x"20080fea814cf80f7c65c68f28fdfdd048ecd6837ac8339f37d31174a2cd9265",
      x"866e9b0bd7d57caf5fc009ddaa92988bbb55049df18d5da49a3284f53c776d57",
      x"648cd331895bbcddea79c8172fb710a5ac1dab52fe3e26e75b2c9415fe57086d",
      x"59187c89d4c92f61c07b3dc2ff61683a0c74e12ecf1e8706c0cbf04d97c6d696",
      x"46d9e893d4d916e02a26ff8affbabc320864624a50398f3d23a3764f80e28cb0",
      x"ac20585b3c546c7428c7ce7d8789754d245f9305578da4f537d5a00ef9792b8b",
      x"99481110467fc7dfd191b1dc55dbdb797bbc35cc1b43487c1a69d49e2a8b5d87",
      x"d2d61e2f35061cdb9a22f83d8bf6c72164e87234ec3bfcd34137e90a0396412a",
      x"dc8328a9f350a60456d957ef0b4f05547cbd9b1a474e28ee4af38c0714013246",
      x"4233e9c3b1c6569521f5585fee27f9826b28a12249ffefebe72283152042e38f",
      x"53ec2c2d79e7d3f19d40d69459bcbed14810fe8ad207357567beab4c283f30ab",
      x"27690734d852037e5b4376a925cb3d67b8a4fcda538befc6c466a5040aaf0398",
      x"cf40cfede591c951f80c2d88860d8e79258439acf601305d0574c6d567f27c22",
      x"684da17eb3b4bee3ccf96bdbfd31badfc37e665a919a6b6a974c1a89ad35c8b6",
      x"c0fcfdb6367021c0751575f172df74b293fa8a4e444f7749a6533103cb22fa91",
      x"43f1a781bb635a24944bb76ecbe3128f9d1f834bc2f29653dbf24a16bb4e7a39",
      x"dcd8580294a09a61621120b9cd1117146afe51ee4f131d8ffad30728114bf224",
      x"1dd3591069c266afe109b9bd11b96d47ea57905d87f6c35c77a1bdbc3d7636a0",
      x"ff80815d283688a09b05261158577eaaa205dc2108f7507bd4a764f21e952dc6",
      x"27d7c48fb6bcd343ee49b5f2e75526fb2cea49ab0e3fe4627467446d0b278e89",
      x"ccbbbba40d3b6b2f41e9568521dde40ee0b00c7eb53f216e2380783cdd6c1e9a",
      x"e359e69129b74c4a6efd0bf969d1bf22cbddd3cb7aecbce532bdd22e9b39a817",
      x"e231e47f70c1cb456f3d0038033f3f75b55f83ca57cad50386ee36583922c812",
      x"98858aca08ec37cf9689f3f5bdac5308cc211f5b9c8e68e6b7739cc6f385b145",
      x"06db9552366de7e6852d9e9f2f2ad4bdea3a221a1c5bee7dad44189cf078105b",
      x"44ed6f92fad538f0c5c1ccbb08b08c454e5b5994dfb5760281828133ea4f3544",
      x"196a87d49d707d0c8898c2b765e9ce086582345a8248209627962c93f14621af",
      x"71f442e85cfc5b1a02c4a036dc0fad0db04e8ee3d5acb63a22fe3e57926475b7",
      x"32c13e5a38c0a07e88afb6d52fe8730d032b850d07e71a36515a18385f22f3c2",
      x"18e848d5679fce47307f8ccca321dd51a23084b17741371284a4ae07946126bc"
    ),
    (
      x"d37b6493d5df44f71d8bf2ab42d40d298c2e39489fc0b7b36947ca6c775f8d78",
      x"5dd3f6b1970e2ac6aafa0b2ff6686753c6fdc744ba9f07f70a4e8df6fa5875a7",
      x"034347841b406e2c90028d4d1e7c64e49e09681aa9969ca0704e66472fa4f47a",
      x"ead01ae9d120cd51af5c2461d899b531eda83386cc631b7ba8ad019e897532fb",
      x"c1d1bb016efc23483f6ae73642afb7b104daa298c2f1fbaf2d247424e10a5622",
      x"f4a596a43d837412978299018ca228df5997cf3ae11411d6873fd5617b1ef87c",
      x"d7f79e9b90ca77fca1fce12a16ceb4024f2df3d0046184b19561c177033584a3",
      x"ce73a014666ebe45c008cbdbc35710eef16149fb321701392af463713bda3b50",
      x"8dc925e0447a855cb3e1ccabaa701e301b8b8db8a7c29ccde5aa36a9dfcc67cd",
      x"fb330355cdce1c56025a66e9869f72f614c0f9106a88aeb589519506a58e0f7e",
      x"f627050d0fffaebb9ebbcb0f5cc80291ff4c59bb48a183a82e7ad90133b07834",
      x"6a0a40361842cd3d25e800cb52a6c059c57d66b1d4a25518fb8e9f73f3750611",
      x"bf4f603206d0749ea771c28c6c93c568d06e6b5204e9e2ba79e9723462303204",
      x"a28789183d9cd61d18f0115702afab022d1fa958fe421c5972b3e913d3f47a6c",
      x"4179cd314088ed27cf3a1dcbeedfe4d133494b0b141ad63d9b3531c8fb49f13d",
      x"3421f0d02c1c9d7824522551041befb57c4bbe2b3f0ed08dcfe6869811c76ea0",
      x"72dcb10142c223c99ee872e482a828896a5fc3653f5605fef737c37a6176ec43",
      x"f36677074c993021b3f06b9320e02cc9f400213953b4b2ac1f26bea86a7f67bf",
      x"4340b84f2ac275599ac121c3a5f1996d6f3e28acabd36daacdbdfa37c0aaae50",
      x"72db244f57e2552aa18e18e39de953176702ee9cec646aebe8b93927b9e389c8",
      x"0b6e616ee32dbf66b34361678c601d5a185233ccd08198ecf9a22c1cb8b87a1e",
      x"0aba93deec9ca1763b9f8700bb04e85e84be212ea1e5acd370fa10eeaf7779a1",
      x"73eee7acf4b766acddae3df46be7bcd4e1a47353f188e81148dff620dcf8863c",
      x"4eb7bfdff2fc21bab25e05224cbf4422545a5ab70cac3210401203fc5d245c56",
      x"3b0ee04c9853dc6a00b11bd26a712c90b7808bf90453ff4d861d8a42afde48d7",
      x"3f84118692f8bec6018ca357f62e5d4894f64c665ca09e9657c284a6064869de",
      x"215c0c89c148fd60bfbdcf1a328feda3f566d8accf370f507610d061ebd587e6",
      x"03f8ea3d53650b483b8e6c742267fa4d5b5d168bb461b795988d3c56a0ed847c",
      x"f12107d46dbad2d6ee6c7168c5d3befe297e28098176d15c9b304171111c0616",
      x"4672a70435a49a4af1155c952d7b1e6b76b949250c5af26e153ca44fa961e485"
    ),
    (
      x"e3f4d16807fc0537fbe5b35a8fbcfe6b2bd2ecd8b1f71bb7e9f56125fde0f30b",
      x"e75a8a04a2d32872e2f27c1a670bf7f0b6bad6db8f875d0fe4c74807fc7b5aad",
      x"549a755d6237948ba6621f2676c337271be46a535e904e92c906c6b4dbcf981b",
      x"d06f7315fbb3f44fedb7389f79891067ee7abcad7fbc87efd3bf395cc5ab46f2",
      x"28d1dcd6ee1b225d19dfb509c8e4eb44ac9de1388ae182b3a881efda154c1fec",
      x"12f910bb17be5ab2601c4819ddd929e68fbc940b650f75f8a6c91326ffd87c77",
      x"c57d150259f7a6c818172b25a47fae6e84dd7bf8dbc8f54bbf9305832ec9d4f1",
      x"b7bdaf7c9c2a40c78a7a7dce7ce964d93ff0f87af1a58c9d3ca7df37c1b27711",
      x"bd160232f5c387b4011ff2c3d4530ee42567fb4b4dab6f016e57f629bd3c0e41",
      x"f752473674c3ed22c9f270c462a2cc2d36c41baa1cf64a46bfd10ed60f37544c",
      x"fdadcb362c6f810e665c141e085fdcf946aff666280a6f41d50f7a093b885751",
      x"ea7a605ff7a5de8f79141d52815bc3f1b8ab7ab3ce046a437a29b284b3c8948a",
      x"84fef99be0bd270114ccd64285af0d7b3d79451c06f8ba230b936a66a4278dc5",
      x"45681defb71a2c1e2df424de6cf3215936e6f503e61180f00da821f249643e4d",
      x"6d6c84eb43caa2a9a2843c1d68e2c6b7b583ce5dded649417d197001a68c303f",
      x"c75e8383790fb0b1415385402bdab7971b7bd2c0dff5b505fb3fd011d156b276",
      x"b1aed9bdac7aa82a251f7f3c7bba251403b9bb62a69f98069e558dd90e33108f",
      x"99ad6a76a288a36e6c5019a17d9b8c9bc2092375f55578636d8c6dc862e6ddf8",
      x"8c9f56571e0a2c36bdba86e7416eae32de3f06393f99744c0161a944c6ccc930",
      x"49ac88cccd18eb4235c58f250a5eea74fa64a184493d6e373ae62c7f958f0e85",
      x"175cae40097ff09a5ff7e4e5158097a0440846b60361ea500688f8ba81101c00",
      x"6e07d5e4d29436a4bf582ee914e0758c0f58ccd38e82dc0d3a1b1e62a72a1389",
      x"05211828c624f7ba7b22d6265f4245681af54284be7ddd6c3a3e5a5a1d1f1855",
      x"309f484af1db0c3f55de6ce2609093ca859d3e13366671ccf26ddf900184ace8",
      x"1219dae1363abd1f7003f14f1442944375c1d741bc793152f1ee1992353a40a1",
      x"6a2034e473a09b1f0149cd36c4ad78de7e3354c3b7e5d726fb1f2f021038f20f",
      x"cbfa8a6c139a2bc3470600842023ed036f02ec1f8854a4b34adbf9e5b567ba8e",
      x"6fabf3c0f04ec49c930349bdfbd5354fc4350c876cf92c49f3ccbf9b93a7c3e8",
      x"1152f14194f0fb2153ba5e84191d81835c8cc65140d915ceb3d7005b3469b02f",
      x"ae846d54cc61b8dfad4f8ef0dee5b96a862e27343635f3a9e83c65c10c35d9eb"
    ),
    (
      x"eb0ed8900747a6db1cd66b490fba5aa6dbe403dda77a74fedc3ca87747104404",
      x"5b6e5e49460f13b49d6ceb53a692d37278e53bca40d4a0587e86f2ee70abbd90",
      x"fe1255cdf5ec137df6005c7cc494baafa11eb5794c94a4a25ac66b1a2c5d8754",
      x"043c7b4a1693a911a2f72f1884fd061ad088bad944e3f2fee2acad5a20839850",
      x"8ffdaab21c7539f935f276fda1b4b191e7d786620f9b06ca7d11adc06edad93a",
      x"a747cce8d6de23c0f26f026b453f0ee5a67f11f1d10021511ff9352d8a56d88b",
      x"2a86b59e94b5ba96aed1051d4649045ab51a19e8e6e806597ef020e57d842ac0",
      x"7451f83cce955d372844d2c9cc351c19798a93cfdba2ec155bcde1d6407b94e0",
      x"dab68cdcf1d8d34c6b281af90df8cf689b21f2a3fe0b03264c80620f5f9ceff3",
      x"fc48a871cd3d35438a8b1782be6f03d8823aca9b865fd0fda05ebd82875cfe2b",
      x"3a05be971e10fafcb69f2e04a41216aa4a44a0089736c9141ccb1e80749f672b",
      x"63521ea864d3f5596f557a410f345e49ac77809757d40447fc1137120e5ca7c5",
      x"d3d14da96b7d9ecc5126f59f9ef7318e5b8fb433a6a77e8f6adc7675513cd942",
      x"e46c81f7b6bfa83f8bc9c00173978cd690beac91b9ee79bf2a6dac2e7922f7a8",
      x"0432721940f3d2ca1d1b44783b91aed2b4087e5217a1801b69d5905da53017ee",
      x"e3fd40fb3e5156ebc76340f174e8ee14b5a0a10f6709548db471b3f35a4d122f",
      x"00802baf197ee8a3f58c8eaf159aa8ec35655e190133578d2bcf0d79c07e4133",
      x"9466dc0874e5042beb7b334acab55d582479c6e52efa4ffb8a55729448d00c23",
      x"5f35a12aefec5725cd68cd5cc5f2b61be4dd1d0951bc550cb75a8705365a0414",
      x"f4ff48c3f51ef7f43c0e7ba1e53300246d0a2b4a15416b663d395af0ddc5413b",
      x"8d76be956b09d98415b9acde317a805c47ce59d01b35a5f359c9d9a30db4f25c",
      x"fdae8371fda7402abc871f043c3055cf1d0a3862ecb1edf384018c68cf31cb06",
      x"bdb4b936db5789c7c96f8308636fb864ae6d79d27620192a3040e1e3bf5bfe84",
      x"086a72b69ce5dbc6ab2ce87f537ff857379d8a8a2c79287611e764e1bfbad375",
      x"5ab37b49a8bbae5851775b6c68e445b38316bae4f101b61263b7b828557700e5",
      x"23e494e7a7ce034f31744d94f50f9181b861f2adccd484049a507c915f74e641",
      x"d41af7bc7f9ec515013f48f07274537ba7dab35d146c1da88da3a1d56cf6576e",
      x"7788d374a5c0bfec239f4f26505f39d4dddddb52e022add66cb01f188d5f37d8",
      x"a48b7904cc58b96f499371151e8da21c243f421a72d9b3bd45e2c44eaff116ed",
      x"f73357ab6415a2c02c602e774a9458037c113d1c670fe433c612c711ade54172"
    ),
    (
      x"c502457bf1962b5c40a5eac705676c93c0c75f7eb25c8924993892b27f64ff41",
      x"f71b2dc1c0d08f7e7558f4b2f47ad544a4610e5c98b84a3a10c5450a96f04443",
      x"ad85368eb06b5fcaecc6287fa4893293e8023fe16422f9cbd1c0d104a422c8ac",
      x"b0c316986d394b5ac656d580e40f9221d2ce8bd9d21ec5ac5cdc48be0fdd430d",
      x"7e92870481bd9c76579f5479a22215356eeac3dd8ccf95fadcbc912b766f3c62",
      x"d6f47a67ca8390f48fe583d67a01a5a8710c024174f77d529b9f914849c64712",
      x"f4cb94de9a02bd338f7eb3b9662a1bfb4b5b94169057332b829bdfd575958329",
      x"fd29b78d38052fea5454e9a10d130f4975ef086d24e5f4e9d7ce8ddd54e5e0fe",
      x"e70195f705e38256aff51058c205510b84beafecb42410bdcef3123cc9e83364",
      x"bdd23cb06b02951169ca4b60c0283536577f081f789057fa0aafae5794053588",
      x"6a65ef6bb92ca64a26d2f022e715a40ba92da67ee03111e506688353db6dfcc0",
      x"b0666c079b33ba6684d19f44909d8070f47875c86f3d7d81b07557f68606b9f4",
      x"497a1b1087a7ab261abd719bc944a8f916e3236005504b71d4a69ec53ddd8162",
      x"cc009193b756caf7faf1ef480321b2ad459f4503789759d88de151eb90d76e43",
      x"9740e224b29a31c5232f19056d05a73579099f57010364d9a9aba41ece0563ac",
      x"385505b08979d9bf1b0458a189d98df6c78dabfc66f30eb08e965df29bf98a5a",
      x"4358c2e03243c13c31c527a84a95e5c8ceb80d246c8b048ac518695d00318b70",
      x"27f9d8da28449d08059a2b4b83e0297fbc40cc5285108604f676689b201a9c01",
      x"542aa67114d89a44d0ee9d9cda664cb5530fb91fadea9f116419063169b573a4",
      x"89f04e95ea05a07f258315a09831718966816655a237e8df17d92734d3fca994",
      x"6d4e7ce524967a3e8c2a7c83eff4653a1a0a80f11ed6eaf784941d2e31834095",
      x"e4e176f9a008b9e2364946573f6b664cbb2710cef9200c93d8fbe99834a1da94",
      x"34161756d06765fa682e6423ce7999b2068cfc1dacf5900f9358388fbe1bac6f",
      x"7f5ce1491df23f383f69a9afa8821fdae8d9b0f7e27d17543dc068ce74f24725",
      x"be0f0be5791af33e027d5d917de1fd52a0b77bc4bca005db9c0c0ebde3966c4b",
      x"a5b4c816adb4a593867f268bf7c57cef47f70474180edccbd8d3bc98e5001e1a",
      x"07160123a62a2346bfed199a1c13c92281448738c874dfd58960524d951bbd20",
      x"0405ce3ef07c27d66beb29731da1a34e58704b879a17102ace2a96c0ec29f4f1",
      x"0a9ee951ab3ac549439e43a645ef7ef33afc2f192930f1a6e57594845df6d5fc",
      x"190713547cd76a7b3b7386c631d3bf6f5e3a9def1fc7ba3cee52f22b9289ae9a"
    ),
    (
      x"c651d6d4ede4d4b621e36b6f305d5d099e585c2eaf44eb897d4cc64e992d11ff",
      x"352bdd5d8688de81fdba1eef6cc89ea07c311a6ef7472de39367ce63e3c70ceb",
      x"3048fa6fc90eacf20b237c1edc46a256e52862173bc6d508bde52f73b5e109f7",
      x"eefe6a34c9c61e78159a739dcd6e6309e48225cc649741b7adcaba5f319c8cbf",
      x"f6dede3e09cb6eb7a97197052e9157079cce19da34757f2d7303f56af6bfcdc6",
      x"71e36680e7730be7d8b0da9556e3baedf6007dce48c45b03285deefa4cc19307",
      x"465a990553c41fe75b1123f75f48f282610fb5ec7461f7a786a5413fc103dcd6",
      x"c545b67d5a7827ced51cdb5745c54e751752d0f51a6dec2a59960ebb7b0dd690",
      x"d5bb544ad39dfe48c75d5564ee23599352a65f5df186a0238f590f10f79ae678",
      x"31778db13dd2b97ba3abd42f16588b4beaedc4dcd33875ea3a4db9a1ce1cecdd",
      x"11e73012c443067f5943120b4b099d2bec0eda30c8e04c8f4ab8a45544aac526",
      x"373a34eb4f7c6d719e170b1fb61a5b2513f7b9d0149836b61c416a17e141910b",
      x"f9d352b9f1f4bea9a1c85cff975b221d43f440099233b882bf7657e72b752100",
      x"f6122ac887710c1787b6a31c602b8f70c544cd03c2694433da729499a5e0e135",
      x"24f4b3e2649532c0bacf66e14650991495591939f8e7228b5bab06e2e481df82",
      x"8014d0b9a5d0d911278f109b5ae6988b4bc089b36a80d5e8a9057a503c112f02",
      x"aea26f0b76e91ab0ff0d44f37b2461b38d2de85d52062420dae43f3359389b57",
      x"37d05bf0e3fbfc63ecc42c8534f85754bf44647af8b9bf407624b1c4edd1a4b4",
      x"50ae726cfb9b66cd8c9828f0c460f0918126275ad1505c5ad18e73356baf6b0c",
      x"70fafca41b17d4f0fd44940081ad62564065f47577f8b83ac02e34d1b6a98966",
      x"e1cc9ff7f0fea2ce7929625ffd36bb167aa8e2b50b5eb1c5380cf82c03f6e198",
      x"ce74afffdd6e43bf6b496d42e251f2c51dfdad13cf3f3f41deec0d870379e1a2",
      x"4e16d4982a1bcbdeaff9f0db42f8747e24366ce658d19a128badd513defc8b19",
      x"0c7a0a0467d21ce5190f566524e95421247522a0581e8bcfb861f42ef8b83848",
      x"7ee73a6c55123f137ea5b9a79242b62f6a8e7adc11f7b744ada695a20687730c",
      x"e2decc8138f9afaeee6934ad5d100f0277c326d501b38fe15e1cf34f56fe4e0a",
      x"4d3247b77c63495199cbea96c9490b48e957a2fd2bece503d71bde5847ad19eb",
      x"c6c40f727acc8604630417436dac23efd243a97fca21b26eb8807053d197e5ab",
      x"8655be9bf666f8523d9404a59eabdabdcbbe5dc753bdf81672ae616c9a37782b",
      x"26a559584d75133ccad0bd38d225854fe0e9f2d7b86d3a612043bc4d7cde1fb4"
    ),
    (
      x"3aea1ce21516fc2d5ed456f0ec485b86d2eb46f81c962fe0e354e04e4da3dcec",
      x"e6d10832148e189d1a26f2d26318069523b462bdc0e4805f0c45d0f89946ae4d",
      x"672cee37800c533dbbecf2f9f531ae0650048c7f4ceb192af5859284bf4b23a8",
      x"3cc72fa82bae02895006994922c2a0bbe6bf9ade6b30f0b53bd83c245b9e09dd",
      x"47d959ce05f6a6e2a9ad23c4c751367ede46634b54f373060f10e01552d40a10",
      x"cf868e35cbbacbd091228e3f9bfd5e044a2d0992d9cddc70be4ef31cfcc72438",
      x"c6a1f5bff613016824945e89a34674b7de1e426b9af51b573cf7992d5d8fcdca",
      x"242a14642c49b37be5443d65c00e7f94c8277958dfd32906a5c664ba992c7fb7",
      x"3af1c6f6045bb6aea792edf53b9297f0fed5a16384ff4af9392b68e5031ea07f",
      x"c6c18b7e7f95a2f0c9f31856d08b9096d8feb9aa42e62c03c77880442d47eaf2",
      x"d8c4cd7c68132f9f3677aa851c8cd510afd429c57e4be0f28d52420cfa75ae79",
      x"153c90b6a1921a668742573d39ca81cb7c30600a0af2a84c8f6ac042e00dc2af",
      x"d72a260ec6b3f915a1f409bbbd3336ba65d169e53cfeffb95f6fdeb9da730224",
      x"fefc76e916249da7118faed8da2e7786a1bc415ad4d79eba9c780862bbece169",
      x"77327cabc72dfbc6d771604722f08a5241c4b2ca192c72f350911a24b843b289",
      x"6611b13f6f261240b75ba9f8acf1705b55eccbe904326e6caa6740f786f7d1ef",
      x"986c879b54ae40c34617ad4cb2f0ee26bd37e5070a136b4ae02a5c76c1fe9527",
      x"533b75c5908baaa1ab063eb570164b97abb5dc271361aa052b627b37211d1d30",
      x"0086c56c05a8f029a456a95ea2f9f5b8d73389e30af94a80b7a2c4df9a246f8f",
      x"f19ea69bde0cb961e6b11f2b79d15a3a9e40d9447f0346023f9bbfd022df0739",
      x"38a9d396b8c52b3ebcc9e050389afeb4bcf860cde934596758b19209165c00e1",
      x"8a484dedd61b858d60cb13a678bda4bb4c826dca2b671da6f415b970c1c39e91",
      x"2edf055af53b77d59709f23228bb36cc475bcccac18e8a691ea2ca84363adf97",
      x"d2c513795dc9c91102228b6dd6777860dd72d526d63ddf1ea856edacd07d7eaf",
      x"4b22f271230882b2ba35ab88fd9d1bbb400251bfc466120b0a65223ef2d2bb57",
      x"263530254098259da490b9600b52a2afa427b20fdacc2ac6c0d594ba320fe4ac",
      x"dd527183b56ca0dd6f7d00a2ec3d22dfb6657584a34d070bf1219e244499459b",
      x"01b546b3893af5b6f004fb77430571be8c68fa44c30b9d684ce7cc85b10f6487",
      x"331a3b777f3133dfaae521c592b0b3c2b8b2cbcc695804d75a33b74260266e49",
      x"c52de8a0524a61dd31ee590bf95d1eef0be50a6d960c5a9f1c5b7027f26a2812"
    ),
    (
      x"7d5a13f66ba46a403731c047e50162a0d45de29119c6cca8c528471d5b8e7be0",
      x"005d153b1455764a4dc7a303f68bbf7b14c6137478ac60555a2cb699177fcdbf",
      x"c9c98c222af5791d8dee23d58fd9134f8c4b1529ba8093e68fe594e876a8050a",
      x"b94930170bc6669cc37f8d4969ba097b9a6f795bf6936c24ccf4db7351e1c22f",
      x"b3bbb8139c64056d440001152c4b1f358d7568aaa42c635574c8bd70fa65063a",
      x"be7433d786e4f2f12290f5ffea7386403fe5411470637a3b6f61da64f4d5a640",
      x"6f9feea8df23f377a920415155a873b0b54ea6cade872bd4dd35cc18fdf25955",
      x"3ca088aec1e04d36caed763bf2a430c55444c9dd8d0d1461b2a564446be27fa7",
      x"7e149aa44e1da5167ffd6e6e7a5de32c264d511c7dc90c45e9366920432c3075",
      x"ed09abf29866c2d0ce7cbd04bd12e2a391f409316c48d47ade083dbc27e577c3",
      x"9ea8cc502309d452a480f9d758e455e4919614839c60394ce11b9d88966ac652",
      x"4d4e1dd456c04174a61574d1ea9d0c805812ce468e16f9035a46d19dd732ddde",
      x"187ce88a7d486ac9b2853680c95e2b66994f5bd938e016d7d14116d931196a77",
      x"292617092eea8b4aec8762f4efd747ab6cac22b375922a3341587f9c987d6ab9",
      x"ee87d0918c5476d80836d4e574a524c9efa8f1d1b703b5b068da6ec43d4bba3b",
      x"dcd8967343d2aeea154128f22d45af284c643bb225bb61dc65409ebad0562abc",
      x"83cea3d69aa179eab0a145184370e1b17aa4730fc577733c520837037af314b0",
      x"a12a5a460a2fc7e5656329fa0e29819f69ce0fb45bf1a88c45736747ba9b1458",
      x"82ce9912cdd9d5be08b7a081b0729326c212e4acaf3e20c08d85ea04bc4f3586",
      x"cf8c434790a6bc75dead8592b29ec5d87ec5bd9268a902a22131edb93355e5b5",
      x"a5926a28281a370499715bec304763474b2e9fd1030e16e668f26265fdfac540",
      x"1d106c4db5bf8a8e6be123d5720cd3573435f9058d8934a9cf12991e286098bd",
      x"4f188de540b44fc147d75f4dfe04863aaab1da222780fa256adbe7cb47485ba2",
      x"51b9ae00521a1ccb4cae0fbe2077fc44c6760dce238b415dc92be01f486ac0c3",
      x"1ba8c251527f1ddc0099ffe78d23904ed9f664ff185116b5f2f87e6186a9d31a",
      x"3b02ec513d0a5352f5d564dd9596724368daa09348944c6f09953bd70dfce54b",
      x"8df5f46328aa0fd924ebea10e2b20c18bee21ead282cc1e9112c73a1b10c8dfb",
      x"37e3963d90c2fcaea7c9f5c3b85fda34dab2159b54e01c882a932fdf807fabfc",
      x"dc9e6fccc98fee322eb307787c6a6da468100df51f5e2e41ea9bfaedda1cd28f",
      x"6bf3f24aba15621eec6dc141f2c854763c415e9e68085c769373270e8c0e1063"
    ),
    (
      x"4a2eaad012a68470483919b73dfbf86c29b9a56248266d107200fdbc185cbac6",
      x"4bc4cc563012317535ef61bfae33dc3687f07dd721341568937ee012aeb09730",
      x"9ca0241e277fb026e2a36edd4ee3626993b7e8b4e1d3da34afa51dfdac4dce9d",
      x"60833b7d1d289f812d3dce212ac692b6511a2f06d196c15998b2764e059a4158",
      x"b148d5a46f691a5aceff548b9f560cc5a3d680b3adfcf48f312439424b66ec14",
      x"e5407c9fe0ff9042915abb3aaa98ee9d7fd82532ab790a433d791c56320d348f",
      x"40f1a841a234681b1edf7eed2e2b3fa032b7b925b816f00a5a51637717368bf3",
      x"a3e0c715fa86805c5b31d2fbd8083866b61acde07f84c20cd62c4f168d7a0f44",
      x"4c598c82a5047b9b5746b790e643c1109f5f8d13ec670e8a894a65c79ef87d1a",
      x"73abf44ca447511acc7e02fae3671eff10badbee6f7672e526dee875ff15f6f4",
      x"056d26d15a3af10577c1e2d781c72500e882702d8c137f6483b4e36439876629",
      x"fb3a7c400436483cf51f84a671c0c120db4d20b43f94a102ec4bf8567036c91a",
      x"9ebab9f8235f3dd6bc9934c3980347359e5f678de52a312e5108e7936ad663f5",
      x"695e45498ac2c32d7576e49fa721b3204e0e8815bdfdf6152c5fdde536d26806",
      x"69545ce62c6a0504ec7e62045b8987fbe46cd4e6ef987d74e025b70d95e72f2a",
      x"170e97f129c86501c1219d4d9338c1191dc618f03af13bbe065ede81d35acfa9",
      x"15f63cd92d6ee6c692574194b9fbe5250a605e1b62c9df7d0be6d097d0532c23",
      x"a4901dc09ac677d6e4cbf9148db9d184e905810ace6d2c8e5b0192f76f8f7e54",
      x"00ef7e06e31ea1cb308ce1c9ec9af23ab47a04db0b5e5163d25c15ced5335737",
      x"415e7b91369d767fd558988455cc6b048d344f37d5b425eafd9f400ab6ac828e",
      x"7d12eeff4b97989cd385062229f5a156b4836a39111fb5c01bc7134cc9d8888b",
      x"230dc3eb83769b8c921799868370f0f75d0631a6dbf28cd1df82d7836d231d35",
      x"36a3327138c7b29336f90b0e8e23deeb33342c8a4594605224f673ddedd7061a",
      x"0d532876f95320e0a09bb035aaa355dd5cbad5d9db52cddfccdd310bd3b2bbcb",
      x"91728758f389387f27cca4f54331ecc12db1b06dc5c345bf6c61612594ddf44f",
      x"bc4155f017f0274f7b3934ab49c9a8ecd46d72ca0cb947ce43f1ef46f09929c2",
      x"e10d9c8eeb3c8ad4d4076fec7614a38a4132fe43484147c1f923117524ef59ea",
      x"d6197227083096fa6819477c75878d51a1d26d0e69787df3545202667e112c82",
      x"1675564ab04c302df9bfb6c251f06834d5b2f183b5790b1f793309db79e86670",
      x"f9e47576060ae0d386704860e74a9c53eaa859e87de53aca579b61dd513faf50"
    ),
    (
      x"2dc4f6b8efcb5851348b4cb88a46c4f05cb69d09d461a6a65858b22290d23314",
      x"a38181097d34e91ef54f3fcb600506abdf3e97a3640aa3746d816f3a6073720f",
      x"0ecdee6548c5bf32c623fd24670353eed1ea39b7b926e9f6f96e72a6efe691fb",
      x"b139ef56ca8696b6f0a9de813eb80d8eda3d7cc3a94af56707509fadf12ccb3a",
      x"c10b89527c7a3b908fb366b2d5da1feba6539c7089305a8df69a57475903a8ef",
      x"e29f6de8b707c9ffa85b4eb945d2c4110fe012e20e78c1d2a88f831945eba6bc",
      x"7976ed02c8bbff9ebbbb0432bf2dd0dd35fcf79d4560c7455ddb8d19827b1292",
      x"a3072208740d45e651dd2142cd3e71a9fac76b480b68f64222046e74676dd4d0",
      x"6b130bd4e816142d210f0049fb8c352af2b1cfef14a1d5dfccee4cc3c0bfc655",
      x"7969bbda86420c3e13e60ba5aa64afe97d9cc7202c8e98a3c5bc6ad85b4c169b",
      x"2c1f7e1b1921d153d4f6923abd5f89ee2fd209242fee8065f9a4781f5ca9cbc0",
      x"2a81cf98d86d3f2e6772a76b4e514a6f0caad6f7e98b6745f5106ba7ea8a3133",
      x"3567168c317e810e971d2dbf9d29fc7a53b659efe11c48f8a95bd16ddadf10e7",
      x"e8c8fd3f8f8ff002673b53968be7cd81af12f51d02221acd41d537fc21643d2a",
      x"ddeebb7557a45fdb3668952db95585f3e81a1378d721230fddf52bf9b8f87ec6",
      x"70d0c490d5c0212df5765f17d4a69e95ee10d0a2f262f1b1f1b82c445355eb05",
      x"c46c9db3bf0811d5e54fd16509848a1e81a3cb32a869f68d6b2ba73bbbdd14df",
      x"e18b4953cca002bf4445d6abb5c5f69f740b36c9bdf5ec1f2db839c577c7ac6c",
      x"5f3c761b21658b28fb33dc81a45e5f97f1826e33e71db2b97795d033404760f6",
      x"3b261bf00fcd31f072353720e30be8f5922f5703d2c34816cb39bce11ec402e0",
      x"f8dadab5a63a32fd048da3afcb35bdd7cbcc25bca7a82e2401261bdfc90e6bde",
      x"0c2eb66d63362df279689d13bbbd8f2520b011deeb74f1a36803cc46759608a0",
      x"8f13a7cd5d38fff0b69fe27b96875958e9f56286cee1d89f4b9aa233bfdb30c2",
      x"9ad01968f38bc6d73dbd6416afb179f6c2d97f62c22004d9719b5bad03c0d654",
      x"8c1bbd4b686395153394544e6dd9c7c7aae9a0233f6931cb6a2857263d97817f",
      x"e0f5a8f3f311c106aa367e32351a0a25975ad431d28a73838ab8a766c3c4fe38",
      x"8ec02b68c69f9a354104315f2d5263777d90da83e80ceb3d64d46edf924218e7",
      x"a7451e15c74ac24115fd3a5d90199901517303c76ecfda75b8e0a92460986068",
      x"6e32c298716634298c19464c006b1acd95a826eb808a004db60e7e873664f53f",
      x"89628ed91bdcc1c80bb0670f11571c14cb3c5eac4439e50eff55faa0fd0305fd"
    ),
    (
      x"ec7d12e5933b7840a42a87c3ba735d38b41b9625bf23c46ddc44cc4746215194",
      x"59fe2b7e489f0db8cfc4aa484cf6c4c984cdf7ae16c74058829f2e95ed67fdd9",
      x"90d83660ee8d8eb95a5dee90d8ea1dc857c41fe7c041dc18f61176edddc8a560",
      x"e2af48576b4e02355f72c56da6e099f4f95c1de9b1e67fc0bbfe796523ff4aec",
      x"ea161a73d0d6b8e0832c08ac10d35595882355904ae1b6310da7ea0276aeb6f8",
      x"7cc69c7466754a672edd64c3079f66ab9abb5dd162f239a642a9909a829e8cdb",
      x"fc0e8dce33ecb32eb0d3768f34e2b2cdebff1056bf396eada07069c57b118853",
      x"8fe9493b291fca294855eea37ae2c0ca2da8b8093fa1b65c887e273415f03623",
      x"08127c394b6d4299037f4d8dcfdd11e62278a9c34d610d042a142836040a97f0",
      x"a6a9c1c21e5e3e87d33babfcfe6a65c09683dcbd50c23031a398326ea1e84359",
      x"a2f402d50e68677a4f3cf67ca43db3c71dd14656e91763f25b89295b4c6d570b",
      x"adb1fce386b26c0de73d00b4196897c7272ab981002d55ccaf5340ce7f1daff8",
      x"08db8d1bcb9114525ee96164bccc479c31208fa8fd4122fce3d6cab5d0980b5b",
      x"be569f87d777a87e61c70b5ac1b44006b8bbc40cc059dfd5c7ceffd7ac1a59ec",
      x"d6e833b8993a39a792e29ee7e07eadfcd68ddd3779cf3131a4406d1d3a8ebcb0",
      x"7a4cba8e5d66a9f55546e224cc8fffef259fdd88a021553a9fbb4b3a70d9bf47",
      x"00c0a71f413a332586e62ff27f3950ffacb027f13fbd2ec69cc87040f560d490",
      x"825b0b0ba2a5e86b629f379c57d95475d8d3d0e8ad61a8c0e8a2b491600732d6",
      x"8d13e7bf66567c36de4919cd7ad75a268a78f2d4a458daadf253e49cc907469d",
      x"fbff251ef61dd549a2ae70f748c456494201ae8d20c1539db6d6201b5aae4373",
      x"f6070e824679865d58d34712d7f3cba8eaf6613c54642243136d41f1e451d1f9",
      x"bc44fe8cd6099f2b5a228e37629c9d514398f5561f38584271645b184ef41cdf",
      x"5784f1ac46fad582f6600f7684ff5b99bc760bd1d9c81a9fe29f6edc49f6fd6a",
      x"69bbc89c24fcf6272023fc36128c1e9f583960185c25e277ef85a48035500ead",
      x"0226ffd6d1ab869cdb7db7a39a86372e7df8da9949156bf2cf0c0e504e3ff039",
      x"37ba61fc24d2f064e4d8924c9f50ce35b147dc174a3d31a26df7f7132776ad24",
      x"e051ff684661f61e87f7e062d7a9a1cf6e83f9863ed46ddaf5e7adbe9382ef22",
      x"84244e905201678639bc61b82b926a76f857f0d87a4ed50b3828cab42a313caf",
      x"69fdc95c7f419e67f07b881eb7fbdb5cf409c4dbb9d6b097625bb159b3f595ec",
      x"fafa2b71a1ec4bd7eba72f1014cf1ae3363fb0fe04f6d8a79dc09a3b632043ff"
    ),
    (
      x"1c605d636f7f9fb74f6a1cf042ba629a909b868c768040b58c7a0531fef6e783",
      x"cd1d8138f8e90173a466032fd61741a7fba892c697f71682234bfaee037e39b9",
      x"2d32b5b1f4279eba36416bab85ce6307d4a0c4fbff8dba96e81a85658f742599",
      x"8d93a9ca0cde12af9cf27ecca0d555fb057caf1dbb68eb6abaec5d49bb7c918e",
      x"db304dc3bcca48c6978979b820b2d5f41ccbe22be80beab51cabf42aa6bd81c8",
      x"a93ccbad1728571077117e5db0ab41d07287c692a9698eeb762f7eb3d4dfa8bf",
      x"961f0ae9b0e3453106521d5bff098948d15e2f6fa126508d6e47f18a33002418",
      x"620568eb7f2ef3b0ae6866f6f019f5346671d8ac77798bf694160a105934b677",
      x"4fbb0c0ee9ac75b110cd3909d5c68c6a4ecf0b08827e74c848267be7ccf9a9df",
      x"02bd94e232997b56ae7cd0bd27b5bd757490ae9b7cee9f1c8efcfc5b6faf8f38",
      x"98ce952d2e2318a916eac2c6275489ab0d1d70e8c5d4fbc95c003bb6052d8cdd",
      x"80e66036aaad4a7dbdbabe52178aa984b6c53c7a8b1d83829b6d5794650ed098",
      x"7ed4e6dc878afc475a387e93e6818f9762e83b4f5fd23d409d2f8fa0960f48a7",
      x"df48fa833ad7de922ec72406724832cb6f95e11c87eb8944205b929c6857f3cf",
      x"d15b157969d722a52731c0ff8e5d1c0436c3e5dd171ce1993fca7f785bf5b4dc",
      x"13cb3d549e2bd46403fd7198a6b469f37627ed19a1fc9ed4deb76b7711d9792f",
      x"ce9f5d029c3503870ae682aa3e1ce8a6c54226b64f178d406b8cb7f4a4b4cf0d",
      x"7dc86ed93df9c2f8a6373fd1c2b0a6e70b9addc83ac0294299f1fb934256eadb",
      x"1d8f114bd934103cf9b3f933aeb07fc38b902c2e8021205fbd9276f9182eed22",
      x"6f4a1c342d0010473cfb7876e00bf78063224cb941e8325d62353c2c581d0cf6",
      x"9b3971de869a90e211b9ee5066031cf606b65f5740aa8d6d0888b83ca9518fbf",
      x"554d6fcb226ff7a8ebf6e5394e8e24d77a9d6c7880f15d78ad6ee33028fe50b8",
      x"7a50ebd5b04533b1501a07f49e84f5beb84185f5f6432a81b471fc177d2facaf",
      x"ac2cbdd3aff6636544dd0a36d16fe080878fc234fc9765beedc54e583b320bfb",
      x"30a560db118ff8bbabd95b6075674ea7f0d1ec89bd714b04a7778ea0799c64a9",
      x"5059c60b5d86dc154bad61ec218b8c80647df8c9da8020615e4e34305edd0e43",
      x"bb6aa72d8d381a028a74687a27eb2862961d1d71035ed66bf13c3aa086aa22a4",
      x"2c0894fcf9723c72427aec9effba77c7a940d609d685b6cfac445ba87d4c8799",
      x"cf439fda896bb48fe424965de2bf9beeb15c645d1d4b5d9d80ea31fc49b44492",
      x"7a557e1f643191ef003126ade4f379ebab5f89d966c750c178199d174ee07957"
    ),
    (
      x"6f5d4d66c5cb92310c5abb9ba4033e1467289951bcee21cd2ab90fddb6f854de",
      x"39ced9bf28a71f469f5d7e3aaa516daafe63d635cc1e62b7dc0e29f739c9158f",
      x"7adb032be8987cc5c16f7d867090502ba0f8edca99bb18c32e619909a2fbba38",
      x"b11807a976d1b8f3324a7628b28b1394d8015a6987f1f97000a2ec4712606bb0",
      x"3d51cc88736e08e43e9df685508d86a48a4b22ec79dbacfead1506b5fa60a4c6",
      x"7f1e623b360de865120b01c3b4c35b1b42b6e59058ea62f43f081fdfb7e82a78",
      x"e7a7910427086e58251c446203e11c58252de165c020cc0684650ec6e1857257",
      x"74d8b27af6f52fbc610cb155cf9ed06950831c023b93351718424eb468fdbde0",
      x"703edc6478268efb8d460acdc544618166122a17c064e88af5c27e5648d06267",
      x"ed41bff018cb694a3766817c19c9c7317d3f6180e98202ec2c96ca54fe854bdc",
      x"f9a78376191c086d46716faab531f9467cabfc89a653b9129679ce031111325a",
      x"8b0648ef4ab775322c07d45e2f2b1790be34558c9839627a12cdb3cf01aaea9a",
      x"e144d540c4114f378b81522c94fc3215e6af38d64a9dd9e76f35a5399072e811",
      x"d08e0b7bd3e30c6189cc073668dd714fb29143ba3f40d8e4d2bfb0d226a75621",
      x"b205aefe3eb08576237386beef6a9bdd627c951aa3ae8734c7d3f0ab04e3c1fa",
      x"50b8893d09ab5b444578e7dd08780350de81873f00865f5f21b29a1289d0df1b",
      x"b59df6889f93eda2855f1e3f3f90dcc50aa26c2208bcf166a06c036503a53c99",
      x"a9ee0029fa61950d1752ff7d81afb4dd03faeaf24244c30364c7825d3284f681",
      x"374ed5c68e718eb175a89cd8f96ce4c1e752f13e3be8ce768e74e3206e3cc4c2",
      x"6397dcb19753e7dbe9c23ed3b2165613ec4fb5fdbe7f54db322e693c7094b012",
      x"7125362054c703dcc392f5b2ff3dcecf2a2c486dc9c27e497d23f641aadc5785",
      x"8d6416e085d955d97ad68d1b46005dedc845350a34e8d86df2bab1e578d960cf",
      x"0946a566589324c4ea8eb4dc1753b578d9d8ea67cdffb1cacb0198ab5c4ddd25",
      x"3dade91b1a68996fc2698e361afa959094d3d5714f496a90f0055e8adb1f42d8",
      x"35cea6ff66bcbdef7e65bce71bf8c45b6ec0ec7e6255481dae0350e126826fdd",
      x"6836062f8d16bca4e10e1ac033133cb2ded76b7bce98a381fcd244790a414ea7",
      x"fe45998cfee4dca10e0ed818cb5c1c0c7d50d7f1afd7e975fc3a190dd93454df",
      x"b4b17dfc6660c7fa477b9f929b729e2f8079f7dca0a86bf85ae5690270e065e8",
      x"a1ec7b3fec07dd77e869f679fb2afd0e844faeef80d4543de7fb259655a30c45",
      x"e4016d3fb9c005d789bfcf5e44921b080c28ccffcc6e4dc9c7ed6c7a3f4a1eeb"
    ),
    (
      x"b6aa1e544ccf088c24e58513470ed56512114de87dd7f3da72b435b2ca5206b7",
      x"08ed01506854def50bab978d2d4f85430472074ee0e34f4ac3c2dd5f06486757",
      x"d641db77065c810c5e6f09873dc1171169cf0dbd67e1281cbda8c6608db5d3e2",
      x"7c2c6e5512a56f36794e42d4f454c23703a557a472d91e5d6f848755797cf154",
      x"da592cd44b1276e32766f84f2b0e9b9fc8eda867ca4c8c029920f4611f0a23e2",
      x"eef8f4fbbea493a298787f7b5ba242eee8325ce06b0843d42858d46b56a4add9",
      x"7bcbc8d6be9f6c2abb269ad26c9cc66fb1a6b5e255b8b20e58f9076b020ca6fd",
      x"cc5eec7cebaae40529020370a7a7100360d92973344fc49a5dfa3e37b6715f31",
      x"68e192de2962167a07a3e4421c56fa7b7666bba79dca9cf86281944be6f47644",
      x"857519c0fd685a9a7b8e4e159d11d082d5006f9c46d27229faf1786a6c1681e4",
      x"a075b72e29bb965a593a69e811b66a5ccc28a67fff3dfdc19ad59ff96397c7bb",
      x"49bc35459bf6dd464dc8a2725542d05ea671d43cb8bd57c464cb227cbe83aded",
      x"c79b351aae912469608f68f3a4db145f8997a9c62611ec2c04d93fa2a3bd48c2",
      x"9db6a1e579f9c2ea88e17b65b273f1eeaf4fd3427e85ebe3c0a7f8c6f51061d1",
      x"339bb0ced85687c445e1c961482e59bd83410f7744029bcfb2700d691a86b2ca",
      x"c370adc99dca09eff0e62774e8824fb62d158509dbaf091bee57bd193f9d4dc7",
      x"e461b93cb6389e494df8ebb42cc51622b496d7ec2fc087f33356f490ef8c2fc2",
      x"7f549cb268d7ab4663635f085515981940709a3ff1cff9c377b38aa433009cdb",
      x"fd721a716a44015a63b657588439b774a285da96a702c0d370371fe9610cc6cc",
      x"384afbad6aaca23469b4205b7ce1c5d6cf7ecd543597f6cdcfd1b59c6cd4d4ad",
      x"6b0530dfc4a3d6e78ef0d3895dfaa224a3f51a9cdd6e013fb8dcdcb09b753e19",
      x"aa030f2a02eed17876c4b483d6b2244faa7704aee563a62d7af27e03d3d78cb9",
      x"a897f88cb31352f485ec351ec6aa166c0d23132570cb4173ad82dca4138942fe",
      x"e60bcc240e1847357ddac6764a4bbc3b1d81ff7a3ed2011f72a8d7adff8146b0",
      x"765497cc0cf1daf6dffaa021f592e4ac58fa90ea6cf4d2002263090294135ab7",
      x"847f4ef55e400519aee9c7f6c6b36a5833262b0508ab6158fa70e2dbde88c727",
      x"b725708b5350311b7c75bd3caaa5a031f96cd5df4968d1a61731fb629f0e33f3",
      x"13de00adef68a23cdab2567329a856bb0471bafa90c7c006f7c499b87b82f59f",
      x"a4ffcc52f5a0a4495c2a3204f76b97152fed8073961f52b5a8dcc52ef8eb55d4",
      x"fb186fa1338cfb09cf97cf06669dddc4e62fb15f9953c521e491f17a69e50590"
    ),
    (
      x"2bf7a28182a56b9909b32d4a90aa3089d93c2dc15a1b86797a6a762780c13978",
      x"adddbe72658bfcd2753cbe4f2cf789b7e2c156d6a48fd602eccde690e7200b20",
      x"0e4af6de14610f4b16b7d7b7aabedc627e1d497d739b65dbcd1c7bebfc0bded2",
      x"22e175731965c47e39dd00ba7b4c417d8e6850a27f66ab0b543f4ab860c090f8",
      x"a566ffe65e1f7a159e46e8320717875531520834c0289cf3ca5529d382b08e58",
      x"1f0a39340a3033a8a2ccde45ec011d0f677d84d2f1f3aadeaa6cdece356d44ca",
      x"7408f78b66a260dc708b3307cfcd6a36444a67953758ed11d8d599f0cf7a33af",
      x"ff6ede2e89932e4122449ebff8d1514086cbe8fd3e34e753feb8fc24053bc82b",
      x"6d494e7a594f4e72192e66dc7dd0dd1f43f97b2351e4c36ed031ce29cceeed0e",
      x"ad4ec5ec627efee859fdb894265769c9c98a7a4879d7cbcecb9ca6001a22ea62",
      x"5eff5f42c4b94850dd4daf898094d959be762751dad1c641c8ca83a83a1523e2",
      x"7291f27446c95fccfa6b5aa86322d893e66505e48f4a3ea19adee5dd4f74af35",
      x"84f3d1a8319e2b4adfce1e9ecfa6c803ba2d46b712428ddcfbfbb61fca78eed9",
      x"96c869e312d7e619e67c34b1201d944eecfed69e818e5077888b81698aa23237",
      x"70db8bd32b191c29cf428d343c031de27294d0a19e794875fcfd0dd13e4b13bb",
      x"63b1fbf81c1ffcc1872a05d5eebbf6922d961a0f318220337d865275559a1fef",
      x"96affc643c2aaee37c966395ae568dedd448a2a27c4075ab2983245d1585df42",
      x"38f91e520d6add1d293625c2597a9605ff4babc3e7b3035f62ab12d5c0aca35c",
      x"8a74085fd2fee480e17cbec041b1ff3ca8fa085e2710f648759b91caaca97cc8",
      x"0b5b156820124226e09e42da612c8940584ac0f8d693d3080984200cb3e6c843",
      x"eec11d7f185508c0e1134c6891cc326e4b5a96a83970c4a64b6b633a35717534",
      x"8bf7fca03c113caad1f58fdbb18a003f51cca999358d5cef1636885c681db54f",
      x"397a6450f8c88eba5e61679aaf74dce5db5ec11fd509ff2fbb6db830d6ef8f8a",
      x"60a4a7c80c3b1b5a6aedeb9a35a6193475a45c7a4e015395193497c49244977b",
      x"4bc7a594dc70295bd5f268dca0ca78fc2db8a188165d3a2f826016f39fe5e681",
      x"c45eced73ca4e32f714d9da961203cf15c0955f7c8fa64a5e0230722a7d233fc",
      x"96059346cf3da4e2af77ac5c79e266982df4a93cf36643e91effedee16677ebc",
      x"cd8c4072d0d559f7e2b3df22fcf28d789679c15b89d7c8ff38219fa02a81c7ae",
      x"5b1ec48c2d01036cffe20f15519e9113011e09a17c8cd672d802d0a9b3fd1ebb",
      x"f99d6e04decdd625840c60d18675296a396018cd2e366c3b0d586adcdd32b8fe"
    ),
    (
      x"6781f76177c212edd36bf642b0ab1e79f031494761e00ea38fe19f8232b1e8b7",
      x"5b23af6b87519eb60db8b8e8258f794445a94194ab8748e1d2c680a3ad368d30",
      x"637da3fd35efa08065368c17aa8098f204384cc699ed8b9aba3911fe7adf5e29",
      x"ea53d67354148edfa08345c5a66248ab085d38e04bcb1c67f0e7976a905b952a",
      x"f7b756506303e58f88210408f53d43b9336b2669256bc4bb7191fa267536856a",
      x"dcbc1f9b4647ac4051e4c5060b69f54c24c2a9c2ff91bd55fdcba5355fd55332",
      x"23e78e55dbc5432076dac433b0705f5cda3a8199be58c6a392803c31633a4e1c",
      x"612305c5d124507b8d4b62d07eadfc5e097591dcb461f316eb396b0ebda6ec51",
      x"c08b27ae149716b26e6207422a7236af30f32bbe26f40c7e002fa29132693c5a",
      x"ab95f54b998b22a5e3f1460cbb8213cf0c7fddbaeccab68bb54d902baea53097",
      x"024f30ff16b53dfd728d9ff178e8f53c578ca1c5eb9b421e965e6de7e7ef8a37",
      x"f845c2a0456e22a308ff4cac1ba9ceb0d7301833a314c621e25e7a3d21d3815a",
      x"0bbd2af3b0419c0d712a3d1119e7f565e10792395323a84119128d868e207eef",
      x"1dd1e6c563a7aca74401b1dc60077f5a6cc0e4a88e17d8e884dd7897ea262fa4",
      x"4b636f63643ae5b98fd4c61d5df08d95886513359b1355729754f05c61c6b40e",
      x"cb895f50416104183c05449d5736996dd589989b6d177663f6dc9f5746ce2f03",
      x"70cea662a3eb1cfe9d436a68c021cbcb1b415373971b2ce03eeffde1aced60dd",
      x"77f045146a225b1f16c9a8220da2ed0505d077c8f4fa1f010aba64b8d9a8f7d0",
      x"d5f5c01063a9f8395c33cf6fc2285a866de5d2a236ae19dd5f8951dc720c83fa",
      x"3b8ebf345e084086cb8b839650d8e74d0eeb2244b4068d7b62a6f4909ac52cde",
      x"795c8105002cacf1c803ab1ec65c0c4dc4ccad86a5e51198ed24387256564eb3",
      x"82b6907068823d6ae17aefc3f3efa7f31622b404542013f03e10275db2c5c0c1",
      x"334c15ba26e5f2f2bd29fa1c1746e46da4465db4c9931e497cc075c274940bce",
      x"8c26508c89e29af21f870c317ebb19e32ac654208164f79474e02ecd241ff8f9",
      x"a846180129771a625f3035396bb993d774db948741c93f4a7ccfa4ef7b0312a2",
      x"211f25313b6bf8f73cf7a796a53f80969d22dbd9e28a31424b60d0aa16ceb9c2",
      x"c930b8c809f336474b63aa549d6be50f0595261a7813c2edb855289c459f114a",
      x"b59d81dd33c943ae75f59a41936f8c95f1eeb10a5438bd2c4aa6fe984435b023",
      x"9131f1a9f136ee0658a171651a2ae96fcace5dd7985bbf00c5089181c1bbc209",
      x"92adcd3bc1a58d0f7c1a661a0ab42c07e60fa44ed011d33918e81d2615f050ae"
    ),
    (
      x"c8a284ead5a44712574f1b6337fc8ba73af146e072d6b880ac64192df77ac9ac",
      x"54756cb93e5b17c3c58dcefa2019d8e59281cc37e434360380181d0f327a8eb4",
      x"891aad9ec5a45ec22b61f02231602b641d1c87414115a798aa3fd046dbb43122",
      x"648cc6f6c98deb82dd35fe04ee634c5f797157c55e8e1d465b7f4073a0812288",
      x"46339921c82e0d86fdb897124c8e1baf95877d062ea448595f422560e41b5086",
      x"5cee0ec6e7f051796e7ed593a834774ee8fb390dbc60e8736116e5e4cb1f3098",
      x"4572cb0d5f49f8330b0e61c3c6b78d8c2a59216f9bfee7ad35b40eef7f0e7262",
      x"d076d7353616ba29a501efce036a61dcdff6a6523bc523bbe2e779e208b5ee26",
      x"296ffb64792b896a29b9e548fb7a441f0088873044edd06b2e9cea1d74cf90f4",
      x"58f85d432a0a14db0336ad6ea36bef8b8f70ba59c2334066b9204fbb35b363f4",
      x"9a6d67146e4882826cb43d2a323c2b2e12c065739f012ff3926a420a95cf0afd",
      x"a7a69e8a9e504db5efa3de0c10c72fc53e82a9a5824e8578324f46f4f6768d08",
      x"4d14f7784939060af57bfbfb7b5a7ed86fdcf756ceb9648d860c85bc5b86e3b9",
      x"9630d3805474edb2af5155c47d7609e40120cc7a1a77a0b7314e5a6a7f5783ac",
      x"39bd3decab32436e942d8b6b2e79520e13c0293ac44e78909a8468d1d495b4e6",
      x"5c43fe9278d9d192dcc0aa68aea09af596452118934391ad6722420a21f3baac",
      x"9405058c43da045ad8e3e823c4ea928f781e7fb03d7fba23b9e91046ceeee035",
      x"c406d22ba4c57e9422e1169e317a1b784050e30811eb23d8a5b86e6f630a1dcd",
      x"2ecde76a98125c19201d760b784622c2dcb7572f5eba61e3410bd19d82860b64",
      x"b9d6bf093e1a9909ac61aa2b33998009db86d750789c46a16af90a0781781c1e",
      x"d443a2aa6b444778ce9dde3b861fd7b3597eb698ddb787398396909173ebb2f1",
      x"6883acc51c684fde348e732c27e0bad64c5ecc92c40b17c157794067e50f50c4",
      x"0938b21b61e6a3651a252e463d75c3f9afd20764cc7bd036d2ad6d2e7558db7c",
      x"2870e9939e824fd7ff8a745a67648d2c1c0a627d838a9f5b3cd17c3f2a8fffa9",
      x"ebe5482a41e5e0e9fd578e68b42dce61c4e478e507a17a07c689beb58af1b860",
      x"b19c3ef582a0640fd92894aba310cab7e06104f7836f25235176dbe47c745b27",
      x"62ca07d2d6ace9813f612b3cf45d8e06442042ee6e7e4122d4ab07d8ebb79f59",
      x"0c17c859b72b2e6bf221d964f6d8eac7f88c063a12c00425589e59297ee24e53",
      x"30cfe7e17e01ac7aac6b6af38bba9260d1bc1eac1c5979c75e5e1190d12e353e",
      x"5da249a28d8253ecebd3af1596fe16c317fae386625f951c80a9403858dd5872"
    ),
    (
      x"89dc4adc8805dc73b0a00dc7998cca509efe6e69ac204a804bd17da244b2e984",
      x"b014a2ec1f7ece5c46758c80b99c4378d603714b3a888c6ff19f462be38ae794",
      x"cdbc39ada0222b74c8a0f840e7c337806757498adfed9eb42d2aed655bbbbc33",
      x"ffdad451eff38993d2bc85766b4bb8e31f153d940bbcfba5daf9a7288390d3c2",
      x"d61e7af440b69a9374c7da70258ae625ea4e9daa24d9e98415382838188e39e6",
      x"762d3bc02e7e5cc25a804a562f86e2b9646b2b11c4fd741a9617fb02624695c2",
      x"550ce4c82636ceb9ec6e390ace37962723e94a130176d2a83073f480b271d3ed",
      x"11256075fe04bbc47f0fa48e49ca81dadcaa85bae0c7765122b7a2bd5b45e21b",
      x"0346ae73073512046e495787be65117d9497c2863726245bf111e7f89c774dc5",
      x"5de6f76a65be545a9014f560ea37914c38a79a07b88fec474780d705520d25d2",
      x"20de125c8e7c605092481249744e5eecfb151ed9953c34405ee52dbc135ad5dc",
      x"06184989e43e109ae9f18d99e6d6988851cb7572e0dc3bccc1cefd1de262a37b",
      x"d651ebed07d55468bdc1f436b2a12ed525d55d391b0da9eb95b32f4071d4a373",
      x"26e307f7a425f831a0b84771a7d47906e03964e4091827169f4e8ab1f6cbb94a",
      x"44f66eba4758133f4b07d8acd96fdcda5a12ef6242c7309a40601e9567456652",
      x"c87ce84e9eae5d28d66930b0df00530b455e373815403e6c724d537614cfd236",
      x"5d8dd264795239ec9126a3ec1408de62f225c69fcc6ca117b071d58dfcc0bcd2",
      x"28a27c61e96f663cdc7d66f92c2fa43c3e493d84e9fa822ab45ee560afd9a7ef",
      x"4abbc2e09eea3e15421af495aa97cc8ed35c41922db3fea96218d5e129ad8cb4",
      x"8f85045e6121f9dbf484b2a722bb2da15fad70cb09e5edecbd7411456006bcca",
      x"9d2aad2ffcb357a6915bd7bfc5e96ec016695f5adbf24dd9a91e6f6166e7fafd",
      x"f2cc0d04725419ff92ec0f56887f2b3638c0fedacbb613a3a11e7b4e48ac2c46",
      x"c5c76d286611763ab8c15a86896a1c51bc4d50712fcc08645ada5711c956305d",
      x"411d310e1c12dff91b408b8b10e263beb8007c28ce2abf19560626fe851d420b",
      x"1ffe7b9be2a88bac66d5f5bda84fe3516efa723f4a76a038d947475b6c88fa16",
      x"0279eb1a8073087e306224f88bd75bd655a2ac7ead3abefe451df9e9f8ad22dc",
      x"5888549e869f138b8e4c38e21d28f91a0f0f1af6b791ddbb83d5807f46ab5c58",
      x"43c27d33546dff13a36c8aa5b61a8663ed3d206b366db88c57fc5a6d48b018e3",
      x"2136056427834faf4f0eec92bf71c0a56c4c38af24391976432d9f633d81b83b",
      x"3399a7b50dee0f16c56002da666c38799f2206b89011b5ac3eef97db29eec73a"
    ),
    (
      x"b7867a6f4a1b65a43d0a59cadba3805a713f35114a83b628cad3cd2450fac414",
      x"c3257cba19c04f2438a9eee89690e6af1bfe779c4f5043949ac3d0bad1e69ff2",
      x"6388caa9c06982c751694c6a14d693a4b5513e4022c97780415b21dbc47d3328",
      x"ee6d177216580c045879dfba73c2c1810574651fb5f6b36427ed693d527c67f0",
      x"5f49cabf15b12f155f433a6592dc5e166539fdafa991eddc255c60bd4605f6fb",
      x"ae43f13a6ca5d59a1b127d06def8597ecbfaef8ef255bc32b9969947a9c838c2",
      x"481f286315563e4f02ee3531e4f6fcc27beec1fe3cfb6245b18db3c64ab39a87",
      x"98f86296d8a4996bc92a36c0609d90922d0adb5d35ac0e3003eaf8200e25b799",
      x"5600f5b58080ea93af08bd8c67442c65b76b11f11a935328c449c9fb49ccb5a6",
      x"60ed538bbcd9023164457f6504d46fceee20d80e73c85223196c77c8d9654d38",
      x"202ef33d04635389b0d4e405e9a54f71a24cd842d5b1b0598b94d28312f2e982",
      x"442863a0c213dbd17e57c5b995ba7addd663daadfd60d869602a9c3ed3b03f3d",
      x"23e953f2fd924800d28998ddc516add76a454de826222b28bd7717bff6cccc25",
      x"007cce6c018ae72d6c3da96ab8d02d342fb667f2cfc1565943810d6e861e9a0c",
      x"d9864b482ba28b036dab673173aadfdc4d0b9c22f5c209e4943b0b0b43e43ebc",
      x"8e254535e93ac688c947074f7772d91d26ec46a6a65856d989511d1a130c5302",
      x"65ed179f9f7f2bd128c7b71ac2aea22d669c8dfe4b53fdc30ef990e87b5c5699",
      x"bc9a389f388f0bfe247e5acc0e796d8f0b147873a9bcf11f6c3ca2ff93adf51a",
      x"0a7f708e81a30a7b1a96640509dc673694c8fc87b5dd2a5fa8aeec78c8334f6a",
      x"cff76ecaa656c3ae823bbc4a4e1766f8391ce3827d817c6ca4924cc856510ce8",
      x"c4b43c1db3656035bf104f4732c8acb8737b15713692c7fe69ecfaff061b45ae",
      x"a4f6a507c98f53b581c69e99004ea5d210da38b2df4184d276c45d6a716cdaa9",
      x"252f4e9aa4cc22e4569cd21f4312f1997604f7aa68038b2484f690f8b5ee42dc",
      x"e63a067a1be9e8fe13480d61d46ffed315e4666584368f50ab7da3e45d71e03f",
      x"b93ff69aa3d0c2390f83c900c8080858c808f4f42c2ec135f38c2e16c1d1f85f",
      x"10f497f5c21aad027544087631002c2586e751a7831ee59f07fb4b9e64829961",
      x"1b3ff8a2c8d9b157a9e908a62998f89544a555df996c314e5d4f02fc26f16391",
      x"eea82614e49961f378848fca7a3076d9abf27e7bc87739b0af7bb7e170e31002",
      x"8a06c4ec686557a626fe1d418264c0f71f7299c28ee5715a4a7093e4be72ad0d",
      x"29222bae9785d33a6e7bf0e0959880ef1ef3efd039e68ee9d545ff8d090c9cf2"
    ),
    (
      x"11c23d3f1e27a16ecc0f53a67b089cd46f28525ae5163e9f25d81e52ee3c6d07",
      x"28fb7bccde838834d3fae08c9696d17a13486f0ba622c0720b6100434c396b27",
      x"d8a6acdcac2ec0319967d3ebfe9c71df302dca570c88dec338f24f053d8cc644",
      x"dbcbded5acde3f45394c444db1bb5967298f9c47fb920714abd380ee8fb42148",
      x"199274bf3adbbd4f2c83cdf61e767ad3ef446c0027822373cd8e732463ceab01",
      x"7edff90b48c0ac999b65618fa8a723b23e4b974d7cef78dd3b99286dc8375034",
      x"65c01e09e4b670dbda9bd1d9dfe3c0534f638ffbbf64a891e1845e093a40b760",
      x"1f044c4ecf5d09f712a67edd99dcf36727884db70524d3f074b26f9c0f12160c",
      x"d50d0d2410206cea546521ac133170b44832ecaaf1ece243fa10a9cf31471a56",
      x"e8db867692dfa6869e131f86e47b4f0246f3101a7609789de848644e1cba11f3",
      x"bcc4b393240bc2891c6cf13457152fadf5877615e3d3985e3ceca21c7fb067f9",
      x"49cbfaefff199dcdd2cb70d0742ecbd06eb7510a6dddefa8fc888b8cc66fd357",
      x"825c6c09dbcf7733aa1adade4dc893a8b5b5afd2a6eb303329e7d702f7e437f5",
      x"c114dc62befcd33cd3fc5582bb045e7262a120ed19ed294226a114e890f608ae",
      x"1f14faaacacd00e2f07761d951258901e5853c6302953227fafe0c24d041be26",
      x"095b0404dadc924c71d03e36b8d41347e456c75869321d127101b37507d1ecf4",
      x"02e00968953a1ac5a565c7e3a41aa68b8f4002b10f85203c01dc5134877b01f5",
      x"cb5a6a0c473188c03bc9c8af072579b983e417b7b5684179b51f218ad269a691",
      x"b694f1ae4ba57b720faa6dff9dd10bcc51a826717f26273f4aed48bdb9ffa6bb",
      x"d0da0dabd92fb00ad93d48ee8b6e916dcc6182adfb35a79a5c31a10cac58f220",
      x"0601cefd0fa112ddd4af0bfc26ddc51a2132b7be9f9e54a9055de120e61e8597",
      x"aca1ff6033e18f797503fa212c3591038185e82bff1f59f5ee54206f5730718b",
      x"829a8602b09122421419b1bc05c29afed306c95957e3e434e9b32be0e8b07165",
      x"e2c66b38b9d8d0e0f606a97d357717debc91b1a7b0eb5f69e6089b238ce6acf2",
      x"37b932c0fecbc5db9fb58af74c156d9e8612acd085ba782cc339867da453a0b4",
      x"5b449645a5dfecabc9a33b2a055917b7b4274126c5a91f2c8694127cf788d3d0",
      x"d595e5e9ac4b0cd5e87412c2c540fa694d1fa0119a17231724328fdae4d4e71d",
      x"1762a53238846f9c05919e33ed16a3dc3798165ab0dc722983fa15c4c228dbcb",
      x"30ac9772e5e6849bed3afbea33c179717cb7b1126367c7d705109e59d76c82cd",
      x"042ba0e8c61959ca9c92dad179b0c7fba50fe6ff197b31b175884eaff513956f"
    ),
    (
      x"85097b398ee412c235133ed7dd1f8922fccd1af55edc6b231c5e7417d75c790d",
      x"a01d931c91cb21faa89d5d2d0e20d116e15fab6e8d35fa07607e70ffa39978ad",
      x"02055b3f188c4b2a8814e54aa9eb694068544b1d26f2c91e81fcc391b29053b2",
      x"4931094e78e19276f43a7852bc21ccb5e47120c8fcba8c5b4e42bcb36b84d33a",
      x"5678bd65f6700a8cbc20462edeb08b026702bbc01b7359f79db055291e02a1f5",
      x"067d840b2d091bb75c5a3b2a90c4cd4b17208e595d15a0c0126197b6a08261b4",
      x"fa8d9a8c0f30d48439d159a3b3c5c2f91af43725eeefbf9902c217625bbb2770",
      x"3eb3be50619518a231b60d6f72397f9fb7bc07b930b4e64433aa0fe856afbd26",
      x"5fe8b47966c5af1aae2c2d6e82edc50e4e2054e8d6a9dfa223c7ab106f90eb00",
      x"a6f3dd5ce70d93cd1fcf7b307b424ff67cf19c33a8e6fad2012eb4bff0007ce3",
      x"953d5edc834921ce23eaf5aef8fbf08b42bfc56ed116e7f2a5cb55f99ccb2d5a",
      x"71adabd78f3879be31db8efa04d2ff5fb7dbecf0fbaeb21395a62536c2010a59",
      x"c3aca96ad7a61636aee88bea498ed9fcfb58b48f18b65c885f4f3e203b7d1985",
      x"04feb9b65d9bb43553b763c86d4ba1a5d62501be520eb6abaafc744f9cec336e",
      x"3e5f26635787c4549161b610f8dd7b38713662dd662956e2c8184cbb2da45272",
      x"8e5572bb621fb03609f20fbb5f78d569e25f96f0e77107b5676570bdc7189632",
      x"5da6206efd1a6fd56877e185791f04a19c6ed21f093e8733a37f82c9d3f4de28",
      x"132fb85471f332ff3994700f271b7caab983f0a0f4c3c365e591cf2c4bba7ac1",
      x"08ae214d96a8037082420bcd3abc357b160bc314e15f67a75874b1039d7f7cef",
      x"0d3a7980012976d811552a59580075ebdaee41dd79194a8b0e1d1f94e1178af5",
      x"5b5a340e61b8a23921f9776fb0443c2f6399b8178fcebc4426935ea287a104e3",
      x"772ffe9639a786c42e4bbd6fee39f7f9a863a7ab52f8f779b6e88ece4d19d339",
      x"9d5ad49bb574e33e3d8ac10b426e56c983e60bf3f3e7786585463b1d18310fff",
      x"cd1163d1e52f54f703e350bad4f41bbc1c807c77f2abc769060ff86782dcb110",
      x"6d57e330bde412acb7beecfe257985ef68c3d261cb10f98129169623193aa43d",
      x"3c4cd740aef6090fb4dc2757eab24e0274242d602fd2c57524ccfa8ab826cd70",
      x"1d61232a1dfc088e2db546fe712ac1dc6b41edc85339afc1ff9bdf1df03df506",
      x"d2d35af9773c6d0f2a6f49016a3a764e99ab9cf3145416ebfa8ab4bdc7cf47fa",
      x"d28987453fe5ccad72f54885bfb139259ac1e9392484e150908df05842d8be6d",
      x"ebde62e2d267a9736a66bb41b6e9a355b24c350606b15d4484632a027785c449"
    ),
    (
      x"3aaceb463e573650c463b8e8c30be0a84a70d72da029ff36bce23ccf5f99838b",
      x"903c2615834016f69de5947c14b8d52c67cd867d0fe5bb1c0955a7ac967005e5",
      x"7fc424313e5e83468c928a222da05ed8dc8f87a66df6199ba5fd428510910f15",
      x"d59cbd504c57c897393a4f6db175d18f3bfb8989da196f47a2c77b7a9912fd88",
      x"a39108b54fafe8e4492759297817bbfa27c21582ccee90d063c82c45dde70554",
      x"d0a41e5b1658137272b9730066a248f09e9a2d02ec781c63d114dcd4505ac836",
      x"7f2774eed3460a83b2375a1dbd083db04ea1a388bd2a76d3d0c313d291296f24",
      x"8233688bee4fefda4dd773630cbe99896a7a374837155cd5de70d9dd08253d95",
      x"bc6a9b5b40096952ac326ced04fd7f92a5efc9903d02b87bd887cfb42297a784",
      x"84e2e8ddbcf0488982ee670fe0b29070eaea23789ec6dbd69ffb7bf8d2dcdb1d",
      x"d7b1f0c7c4b998fa2629bd91220237b778be5d3d2063f8d60bdb5dd5a30e9e31",
      x"c3a3efd1e2653497f475e471cf92405fe91c976041529c80046b5e8fada8ae6b",
      x"726fe65371369250168f49f7f5dfd42511c7b37a78f2e3e348bfb17562d6953d",
      x"b61d108a339074c19308430a621bf967151eb5545d079c6ca5e82f4b76b3db2a",
      x"f3602db698ccef01551648e0d403298142fa125e5d6c5864bdae89d1a49b4b74",
      x"0aeeb9ad5349f63e3a88c49a1767c949ed08299d29e298dbc17309f862030ff4",
      x"f5ddedc3276d223ba6daf5cb4c7b5f5e42912d78e91092451ca8f7cf3069a4f6",
      x"0ec76a64de33cd7fd05032df3f4334c0de86c8c93d64ecef72887c65f23d789c",
      x"92b5b5a6030cbc4bd9b92338bd5a6aa365f0cbe225d120807222d51306123acc",
      x"1717b6d4dcbb362eef90dcd16a6f2f0659f12a804a56e95413cb18f9c859446c",
      x"6d03725a80c25b7a072618af737325ba2c84d7039fc1550d70181a60cca68dcd",
      x"d5609abbbf0d179e169b26e9dbfdc22e43f851470fe2717c5e9b072a284e8712",
      x"06a985310a651d1f20b0c8438227a2f714db9e180b0a54aeb2b59b5cb975373b",
      x"608114390003f1cd55e7bb8e254532dcdd1ec1a7513cf040a2533c5da588d4e3",
      x"d1bfd4f515ae275ea357d8b9ffba36f48a174a28461fc42eea9467067dee9c18",
      x"e583a5915056fb65d1e56d2ee924ccbebefeb4922526cca2db42e29bcf216f7a",
      x"9f07d1a7ba62a52f35a772dd6b00423ced6f765c96a678c2f1a0c39140012020",
      x"feb88b223737fbac7aa51c493a2cf2ee884cc9c0203396798636df11ebb26356",
      x"11ec68dd055257f2369db33d07e79a5900f3d9d796f88e1db11477b3d71d03c4",
      x"d813c1cfeae2140bca49a0673c9392ac6d503da81ba6beba21ce40105ba6ff0b"
    ),
    (
      x"e468b686807c8becfbd775014ca0c91cbb10a6d172a5b4e8027a8434756dc940",
      x"47ac63834e70a842300ca12663a66cbc8494d9711efa8fe71566ac2237fea697",
      x"13d88732e734d9d017f7b95436d9bb372840ff93bee6c2e360dadff156f30fa8",
      x"0adafef1cd07db7816f8ded559d4475ed66f0d0b28815bf6493a2daff4992539",
      x"7c842539e2d383ec652091959dd6c245e99b4195c830f3041f25db5f916eccd2",
      x"1741ca93239e4a24bf4cd5995efc09474099c241ddd5833771c66ce835ec9801",
      x"6e3e975aaf7eddc9ceb1c0425174e716f290a5ea982e6dadb31ea8669fb081f9",
      x"1da9c41c007114f1627f887876b566b70bbc7abb4229f0c88c8ab53f13e71c02",
      x"74f0236fd49305eba3f4d9a5b8c2d257ee007978938caeea5a05457f7d737244",
      x"fa713ef2362d7df5dc14b406d4fc04f23634cf272a0d6afe3a8bcc9b38ea1930",
      x"7cdbce69cb892f19e17bc1f04a50be66a91b90681391a296dad35578cf61295a",
      x"57817c0b4ec12d9b5843d4858525716b89844fc7b59aff17ff84fd1e2b648586",
      x"a63d63bafaab8a0d62bbe4193dfb0297734f09ee5a694634a5cd71b11e18b6ab",
      x"7b5c3d8cef86ab4990315172eeb60437586bc5ebdceedf1acd8e2baab7b23ff5",
      x"608d18c89098984cd07425a17df2c8dacc12b6c3de22b5d5ce11f2c4fe54125a",
      x"a30c7638dca370afe5310d62e388684e11a1e7ea41c398640a8c7bfb7004c22d",
      x"2132ac031da791af3b48bc5330260c968b18bbd71d392f9f452ce3d6edca3d2d",
      x"3add4597e0a0b70186d13b206a048444b5a37dcd8748727728a74b924c7b5be5",
      x"fa380552b8b9fd5931937e3e786f8354bb2bf5883a36351f70904f351573c9e0",
      x"3d1f0703c951bf4211b38eee264232f7d47d56deaf6610ebe84d8677d771f4c7",
      x"0140d8a4354eabae18a728fbecf4354d7d54433bd3c6912c3ee7889e78407259",
      x"45a72459a982b5c27aeb71df7b88615547ba6d26a3e82292be6fb992e2a508df",
      x"2062b433675195f2fe4e0a622e0786a92f33abda565f17a66b876761c83f9df4",
      x"61fdcb88218c116dc30f75ee147d24f355c60659101fa90dcc78bbf5caca822d",
      x"a6299ca11b5d38d5f096619fad341f56781e43f4ca6a6074168c9cea064e2bb1",
      x"9a50b60e73283b4e41d07c69466ff70b812acfbc7519ea860f4aff99c1ae6ea4",
      x"4d36b55e0a889f1821542260b9e63c7fef3dd2eb68d505b8e0de2482c4948fcb",
      x"de2a788672d7aadfdbdb6bca0224f3a6e1b543313d14025d80bbe54b521b3cd2",
      x"86938d1a74920f9457626ccf80da3281a079983bca66c03260e310a216eddbec",
      x"a77361cc2d0a6b19adb585d455953a11e0e44c42802b1696b763064f78e5e61a"
    ),
    (
      x"1d702201d266e371958f21723ed5fa5886cc7c68619a874ce7a66dbf6e0881b8",
      x"661a94c39dcd56d88b140758abff570c002db9ee03c46b3bb6b531d686347a51",
      x"6c94c65e045b9bc6737a1a10c97038275463b62832275f50f4cea186beee4fa8",
      x"0478f8d61858a5f482abc98ddd0ba055f18d3d21ad6333803100d85bed7e6ba4",
      x"f968d91a048ba8e515a68ee459ef12f93d2c3a9ffab7fa0cfb6199840ae202e2",
      x"9ce3a27578f98cc8e20d0948d49d4e023ad697bec1b41b7a3188977e5926d8fe",
      x"775d514f0e0b12abea071fd5515c7f680c0577bcbf73792da1df93a74cacbc99",
      x"bb7aa4a7fb049c3bdf82ad304f7376f3d6a841d36e766ddb8a876f259648cc64",
      x"a4cdd8f13de2b733c7d6f320a314a2619fdff5f21f95116f0e98ccccf60df303",
      x"4a62901ce57a914ce7960b59ea771664b5a4c306a9661d612eaea5d19798d7e1",
      x"b1177895d1814022900c254eb344e3b1f8aadf7931cb2d092ccce3e583369154",
      x"1c2561e85e660147ad55bf9b7d4e380913142e782bacccd91d6268bc3651a1eb",
      x"4abd068b2c1e9a283ae74127acad28dd5389f351c0079034945afd0b85523c3d",
      x"0d197da5f5ac4f8f599f0ecb8f2c46d61a5898db294554091bebe0121b12b2f8",
      x"a1227d2e52ef2d7d77eeb4576ea8eb379e293ef34be2a9b48ffd322876ba7e12",
      x"d40d634db0e6a99b0b0a8e1170a8ab9d9a8fcd18f57f3341a0ef413c391aa5fe",
      x"3e21d340d1f263326c223715424fe6c7767201117b36eea728a529adee423059",
      x"57ecdadc551edaba2a53c41ff05c9cac64281a1fe147acd30929ad316ba90e8c",
      x"f716ec66cf96d180bb76ecf677731099da316a6ae99ff4e44b50dba59fbe3803",
      x"44812823db5d42682539a1c46c34e844c7cfc95920514d08ee060f839b1d0e4b",
      x"1be9bc3f21639f8a8a21d5ba8210d30773932fc44576aef6438cc48662d688d1",
      x"05dc866d7f637ca1e2a947135ca4eb1df57b868b4846ad52ef452bd91f296216",
      x"d74b7c4f5a71b7d27b38ff0a8e39dff2550ae661890633e3d9000e4dbdc8ea17",
      x"05d2ef76732a17c7f4896a21a5dc8a5b682962d490df8fb0e7b9fb3b8ecffe3f",
      x"852004469e5bff0e4c3b705152cbb433403ad58d645a60066d138faf927255c7",
      x"e23f8272b766e68c8e31410e4c8aa2967911138c7da28e650d6d0216309d8d7d",
      x"461e4a9bb1360a1d1669d26660e2f3ab588699c0bfbff4e0f8c1af4cd8e30d1d",
      x"1107e348e8e274d3640c0a9d635f1109c20258dc7902e31b9cacff7672c7432f",
      x"eb68d3837b28ea63ea553c1bef211ac754f3ed080492d682baa85b01db33674f",
      x"e26339bce1d04d01dd9aa10bed251b3b59f5d383c80583a11ec4898d94821344"
    )
  );

  constant ZR : T_NN_MATRIX := (
      x"8eb5f9ddefe1974c21c255023ff07427bfd2010bba4225b16070ad1b9818ff0a",
      x"fb8432ae9cff796843161cba41b38647c014ad82b55637641c571b45a848dfb5",
      x"6fe002827d4b89e9c162b08b8854cda982ccc89743fcfe2a0aab474ecfec7c11",
      x"bbe98641a66735d82ab3ee8e020985a435091e6bc2117abaa9a462d0f420ccd2",
      x"30be63aa4d97226371fcf7c3a1ff80803a1eb049960a2054d75714a9a01fc6c4",
      x"82c6abb46cce93e3eae50f87a3dc0072a3142aebc96a83e027b34436257745d6",
      x"8677064e96d7b851fdde9f4afa5217d1fc4b5a4882d513431896418b61568fc5",
      x"51c457e45a54b3d7e2813b8ff23df05e6322e93599ac08166ad63e0b3d9cb110",
      x"30bd0a3a6056f281b8b61789729a62cb7364c8fad6b229dccfdfb544a462ad50",
      x"c7c16c01fb84f65e1c26da0df4b13499604d2a1316a5c68342df8a413f85fa1c",
      x"fce5fbd6af44ce90d6548b5d01e955bffc8910ac88dedaf991a9fa4d9da78a98",
      x"61c72661201277aabba804701eb54d08c672bc532f15483de74573db4c062dae",
      x"4d515b661e9deeb1ca8a9d9b05524e71a9ddce8cc1e54d1133fc36a3ac6cc248",
      x"3fcebc9d020506753a8046914f5d3c702508939d3e530d2406ea9a512700dd75",
      x"aea968a3cbb115a5faa4aa649f53709a909386fa98dd2fc468c3fb0bc82e265d",
      x"71c0d99a2910fc5ff860584398360f24ac2dc112aa55ba619402db0f4b063811",
      x"8925ee24f2364094bea37d1b27917c403859c3b355f4f82da1e6eb674f92f74d",
      x"4a2b28fe52908a1653d220258a9c4b044055e459fa2821d2648720d8a9e3d23a",
      x"c90325bac66952a00a0c2f69b2fbe26ecc083c14932b9a87471a97d99f7a2854",
      x"2fd7a7894272c0fd99b5f9ef56f82d1f799f8197ab12a5f9797735ca04c6ce5e",
      x"93c67375d6ef87f455e499b0db6f9bc69984228eee2218af5b9f22bc5c673f36",
      x"c39d992b847a0a629aa7a9a6aa29f6914ffea2dd0a34c22b4224c4d84dbb3066",
      x"dc16a6b0c0ad4e2ded9b6d48ec806978529a1fb80dc23673d1f8848a881041d2",
      x"474495e84f1c3a22225a52ababfa21da7d133cd0d52cdae69b407a916b4c34f9",
      x"18eab6a276a5befeff863392a6fcf08458694175c862cb9c4364908e8818f1a7",
      x"a78472cfc2441158a6a73c050713c85a43bf7929648cfcf0ac24b1798f71bc43",
      x"31c760b7abab11d1ae1e71505753a27fbd729f61b78583f60ce5ff1720fc01f4",
      x"bb304157f980cf2b41537ba09e1348f21bfd4cf8ebb41d20608f083e435ebe64",
      x"33d3facd94b9d0162c87473a7ceb91a29c6882a3c5909a3f0481bb3988b2ab33",
      x"beb081644db71b7cd952b3ffb8c84f2c5ee63f98a613f5511957fd9874da89c8",
      x"a4fae5610fb8c57d361b5133633529fbe7b84a30eee2e9b4326d8ad65c531aa1",
      x"66ef969a06a6a0a8b2bcdf9871e17a876daf4faab3cd5caeab1e0b4531966369",
      x"0725521795411c3ed9c23f8e0edd8430fc5892c67323bf35a9fcf3672dc88e95",
      x"eb1256e8676aa708ea201432fd77ef777d32e6784c54299f948cdef3365bfc2d",
      x"2ef5b89543cfe97d3f538e2dc22385aeb5fa9f57f10bd9fdd4527302bb6ee670",
      x"da030b6e6a8f61c6f10ea84089db83cd796becb7b42f731a8c425c393da15b60",
      x"bcfac35839605ba620d77fdd2e0da9762581469de10ace19fb16e0e8e434d4d4",
      x"15cc9a0eb9882e748cef67eeda81bd0d535bcdb6e756f85bef776b891a8258b6",
      x"5f42dc8370c34278c1bd08b0aa358eadf1e14019a7cb053ff43ea54fd3675480",
      x"dd83de7b87eab63efd5614e054e23407997b98fc99a95568e14fdc729a1173fd",
      x"352e83117ff2ef321045317ccf8e48043f1049769079e78e8223ab7cd10168f5",
      x"4677753ea905ca7a8e3c93e2c964de6bea2ab513d7b899f39c502ac9bf3769b7",
      x"365c40b4ce7b80f35b74c8f0b7b056d2ba0c7bf766e848f1938c182ce4400a7c",
      x"48686c30602922e539484c45807aa93034c4810a50000592fe264d590b7380a3",
      x"fb0a22a513ea98778c552d82dd55832d40361fc7f8b389d44fee901f658bebd6",
      x"097f50afa57560d2dbac05f19a05acff26c69340a4bac3ac8632c05d35fbfe10",
      x"ccd200617232178f7c6a1f6ccaab7ea4e9d6e94fe7c92b16c4f1eaa1e2166a10",
      x"cee298cb460d0febe25eb85b51bf46a3701dd2d406f06b8cbe3f604e4a6a91db",
      x"0744411358e16b04e2a0fbf0968190133b0080980847f9502607c723db900660",
      x"df18a6ba512ce0bf2d1f0d3b223cd390eba7dd48dea9aa2e802a6eb28efb6583",
      x"3dd6a9c474af998b57dec4c212f757f0541f1898137fe752e27ed55797f51a2d",
      x"5251015e3667fd2661048cce9ce09163a656f2d1e07b33e45ecf15bea9e1e506",
      x"e491d6a51165797fe5fd57addc61d394cfa09a46216d1506563d5b845ba80365",
      x"3036b9d1563d659a79623656cbf0be53f2c8eff348bfe16cfb0cfcbaa73a3d4a",
      x"134b9584915167c363d0b77a448744d5ac9e0b12fab665fd9ea7abdf72f0120c",
      x"660b153964621912d60124088ad15ad145b445cc89b02db6836a08627f8fc796",
      x"495dd0e376ab33fbacbd4c589a04dcb6341a54492102c792b655f94aa6e375be",
      x"d24e1902ddf57ee56f95f9f1c944ab2f9b22603976068b930b82f3d0c7bb3c96",
      x"83318252ab533dd124f9b9e6679d48e63bf07d31c9798a25b302dcffecbd8a07",
      x"42eadd002a737371a17c7e247def1ffc64aae8c6b93909018cd9dadc65c58583",
      x"0366466ea2a70bf330be9f482be58c76f1b256750bc4a05a440159dad3e8f26c",
      x"08a4480e07322c7ef5d6470d08f3c342354964f97407de92ccc0636fbfe13536",
      x"410e1654cbcc497d5e3340007e94e660acd10b04b835fc1eb523d3118d20d0f6",
      x"04a765635525eb2d5c86ff782bf1b1f72b5a93c44ac7a0648c0cc2e2962213d9",
      x"130b7b08225f72c24a949e2f9fd9b8359d5679b0c8ec7832deea4dc766bda848",
      x"df282c0c1a9eb13fe18cd745c134a09af548c83b6203734245c6ea020065083b",
      x"e0eed8ea267067ab98cc406bbaadda0ea88c425dafe94800deacdca630ef974a",
      x"c2346b55c784324677d86fdf109e9f85f458e0229e249d3205fdb406de2f8fe3",
      x"358e0ba126e44eb0026cf65dd6d15410a9f0b503a26b06b4995f12a1f9b8a5e5",
      x"04ff4c76eeaff49a6f2f8168ecc6105de041524f215eefc1b919a8282a99b33e",
      x"a49a096d19dfefc83fd66a8103b9278512a7d8cf8d63fd2692d43bc5ac94d0d8",
      x"5b8026c53f3afe698fccd0bd5081d4f3b51e868c09af4dd1beb39973e4bc2083",
      x"320a55de5c40e3e2ad1a7a4967d2feb0721b825fe752d486d5be831895ad62db",
      x"0d015035566b728d474c8a3d628f9dd8e7c00d337007937adceb53b0052ff528",
      x"db349af601067306e8c26bb89b98da7c70519494e1382c4b415d5a2c50410d02",
      x"4c848a8bccc118d4e4d8f8c03cb179d96655751df5651003dbe97311ca826676",
      x"8499eb08d0409063b8bfbe19ad3f24504c8471018ece24659040be2674ea5df2",
      x"5068d55988c6f35f33f8a1d7fe72d330f4ec61369ae85d5882f61dc78ead91a5",
      x"ed05e58b7fe327dd03d33373202a514b4dab4db5bc64fe88ffcbec04035a0179",
      x"0073c58ecb9a230e528255a70504026edf8c8d0a5118b5d70daa4a7a0a16b364",
      x"544515da5563d84b0675dc0d9d7abe82b10f061bf1c8abc3630d14b1eb6ae96e",
      x"188fbd32c05b31852000f8bb8a0861db32254617abf1400c286df8bd85b844a4",
      x"e35529e1153190becefa93b20fe8c0ee1b67e31e0583f11ec51b80d86eac611a",
      x"2de91fe97ce7d51a755b6f507b6482bae1911875eb80ee87daf39148205165dd",
      x"5cb7c2b274395ad3eecc1e836476ea643cee802af2c50d574f04cc16fef88dfa",
      x"85d49b15b3e020a2c79a15cd9a3c0f100c3097e552725e80ea6564b9050fc94e",
      x"a74b9af74f0f98f4546b1de96b632545073a4d91aef4a16f586046a785828f2d",
      x"87e5f5394c78354728ac5c5f2e33057ed961addc14883acf85370ae6d013194d",
      x"9e01f74a135f874c51d1702f95e40fb9c5d9334e20831a652ef89187c282e24b",
      x"92ffb578db76ccefdb3782733dbfee9d3ceeeb01dccb39220f32542a197447c3",
      x"44064362b80ea10942bb96735bd18fd910727f1420c3d0eea9a9062b6cd71fc2",
      x"5a61a448e68053bb99646bffef6278b8ba8a311b0fdc49f956cb00096db8a8f9",
      x"cbbba3e9fca5f6717214a9e99c847919fa6f6fb65c31b61d43c0309b5a368ef0",
      x"09694124a26d4d34675f3f2bac2d974db86ca2a34bb567b7ecedf7c30504f72d",
      x"7070a497f134f24a0d57b302122ad5404be29d4fe5845d3d152eb895044e2e86",
      x"4a96273019fb9417abeefc6cad7d9dd89d47e0c618460845799ebd8072e58e21",
      x"6d3f399ace6c111f7d7e98723b237bb7784aa47e66d34cf48cdb52fb76137507",
      x"365fe160161e446547330e7330b795c7d5f89639dafb927da49113bf2d22e72f",
      x"68d4ac37c4c47a268e0cb10d71c15dc2e8b2243d4bc1fb61497a2ff8880afa15",
      x"4e650deed3d4ee0384dd78b09f306f8d02aa75cacddf2d7927909de83bf6b130",
      x"87f89fc412f4238ae3fa1b11211f228e98a4952b7330e86343c3fc231e1be3e6",
      x"d56fae5b5f760c79f4c00dc3c1f339dc50e0d0d0ed1a150375290f2415ef03c9",
      x"b369e8b05baf7da974a4fcd70844609128cabce9c577a40b1bde91c13a35050b",
      x"f52b97fe997b5cd272ef9b735765fa8c8c79af65e5b4b46a9092128b741a1523",
      x"6435a6572a2a8eb970ac078c05c2b9b4eecce7a02733ef01c485b3a8b404f959",
      x"6dd99ed16b1db66b449a3d4e3143240c3c52c81bbd695d9823d45851239b70d1",
      x"471e0db2644b245bfe5453a72646a835c2949c6d55f341929e22328bd9905077",
      x"09aeb8e2c854eb5fcf62079367efc20c3633cef8075a1ac41f512e8db2f12739",
      x"c41fc4f9a100fef88ddf5582131d44c7db3c0e4d80433c964d60dd8f2b1ebba4",
      x"e80c9643664fbe87d9fbb6ce7b2ac7a91329bf8eab79e548d6f1b776719b4413",
      x"8de3cabb89c3b7e789e68c3d4b2d2db00b2dda239faac964930ea3ea2c32e259",
      x"0ab0d57306384248c1adb1bc3a55c52d67f4f9e209c707854777299859f67b56",
      x"0aa86c6e305895a78e31ba700c0675fe6445a439d8cb5d100ad10a025b04f924",
      x"c9d3896c821ba06d62cfb6cbaa1f62e728877b33204462825a949a47865aa2f4",
      x"191f31d7dfde4aed47da2bee85558ec335f43b1585d4c1f4a520c4c21757130a",
      x"91658646f713b42298d3fc270afe7d58bb94bd380344d277cd92825227eea14f",
      x"7e9d079cd944726d2fe403c52638ce3e3a03b19273e73f0a882c665d60601224",
      x"223a729ac4e0e6a42c4ac914640477b2ae1479e4cbacf079ce921adc2fe34280",
      x"6afa7f1973d9a23654e5be8e14fa30905902152064d1602ba519bba93b1c961e",
      x"3e765275453d92a691ce98de5b2201a5fc4b69f0867332ea4112a71a4f98f75f",
      x"cc4db151e3e5dcdbf635c72dda523241fc4fc890633c6346b5c8f5215b9b9700",
      x"793f66dc55fa65b1f67d28b5a06e040b3a8badbaf083e36fc5bda7b4d6ff07ea",
      x"446f29ebd9cf9a2ffa6d340cf86dc12689a4060a0f0fd7a2abaa9148b1da071f",
      x"7628cbd60d887e48b1e0df20001ae293c4d667b65c0c960450d18eca6a332564",
      x"43e3ebe72deb333708c42087e4a86c92990323ea6b911f85e8edbcff82dcd355",
      x"be3ed9e5ddc7c623737cafa26a32c24fa39d1bf071ab693ef5654c0d3406b310",
      x"87d19a98dbdd2c59b417ef60123f87913973ddfc8bb66c43d7550c764ee16407",
      x"5ad2e039a048cdc9b122302cb7d9ae696ec8fb5d383e14e237838c820dbabe29",
      x"5444197f1cef65c09a9020cc8c36742a5a1c79498bb5361cd7f62525c5d367a3",
      x"7b90f91832b40bd231267e093d8d88af444a366cd5dc0763866f599edfa9160b",
      x"9bfb1e23552320654dfbb9b43ad636316d9c42f674d74c1798d1769657474e42",
      x"5b61fc1f96add70e41348b8ac45fb004da0338f3714828aa73799711773b2c6e",
      x"0fbac216286fa06307934ac6740e6503312f4c8e1802aa10a72ba2f3818aaf34",
      x"e7372a64c711776afe702503878a1bc31f9492f09ef2eb362fec2a22d1c5891e",
      x"9071b6c82aaae908fa8e17f998de64ce62a8987849162292898b60ca170e03db",
      x"38975255613a127a9713cff2f23f250eb9038b573ef28f17401ed9edbde1b5d0",
      x"495dad951dd1b8027a745ff64de244f28419cbbb871713f440c4ea942dc116e8",
      x"5268fb2134f813857373c6464737464e2c6bb83a30d138ccc96acbee7b30fb7c",
      x"3ebc9799b6a9c907c7c4cf4048965ee9bebb515c039cda241e7592dec44aebe3",
      x"9a5fd1c24299286b1fb86f381b51da73f1ecf0e01cb18b793c79f71589c500a5",
      x"05d648f5cf7ebfdaa0c37c0dfee66e434f701f285afbacf9058dc1618c252b04",
      x"75c965cb4b4f51103e2a25286e57680b7d49dfa3001a9c25d36dbe88b9cdac2e",
      x"b332f27b7087d0c4ed36fffcf526bb90a5e783bbcac5da527199de6b4de81af7",
      x"e5a3d5811b0b505ffa6d8a0efef7d2f6404d2cee92416c0cbd651be3860bacbf",
      x"55b39491f2afc8324ed2c2c1be2c5891812e497b72403688a6d20e29856f80bc",
      x"d40f1dcfe629d4829887bdd95a434891ab4ec20e7ecbc7085852f8a3651141a5",
      x"1c6f176a26e00a5d7ec74dd74d38e55ea5a1bc6405d8dbf1c3032495b397fe2b",
      x"79290007e59fbb4a684c9f814708941da0afab5fe6545c8de197618986f1bf29",
      x"1bc4b1b9a60432bdb1a851d1906e1c56609dcec322fcda579e75f28f6cebbe3f",
      x"f587704d3d8168bbd5eef27b7c2061e5f4b9aad9903e7a26417f9369cb61a987",
      x"1eac4fafaf22577397e721f0415feec89e902d067f07930c646a40e34750d8fe",
      x"12cfc6c659c82768e3357c6e40daa7ea3db37872889341249674914162725d53",
      x"67c9766bc925362e4a21e25239bac204e00452cf62a6ca1e46f9124f1a8e8775",
      x"e5d18c7c25cf5dd71e812ce9ac4704b4f0785843c3f93e850319134d73b9ebff",
      x"d0487f3af3070f924f14f32ce0f47466f272050c99809edeb7578d01ed1fa117",
      x"3a81f7a9e2597c38a6758442ba49ee90a63aea1f9a84d200aa0e7c8fce7d29e4",
      x"ddf5f0816e2d6ca75a27030e66c6ae701ae9fd754eaaf20f839779e58f43ba51",
      x"83c0ae90c4a1b05ae66d94b56c71ff730d8f798b2f46220947f1836939275ccd",
      x"e66607d18afde80ffeba6edec4ee094275e2c3fb0424cbd9f29e75c0ee722626",
      x"e1bdc8c0ef2ced28fb8b604ec6d659c5854f894d5a20130e6ba3cadf1db504e7",
      x"9cad0916156732719e8bf607f8d80656dc5769677e8d613cb545ff5e12dd40c9",
      x"98bbb1920f90fa987851cfb8d0a1c225e2b23445f6a705c818fbe36a8bd9b31a",
      x"a59f8f0fde7628f428fa23af61bb07822135c313647634b35737e27bf53cb559",
      x"9cd190f4b17914122e7cd8a1b69c7ae7cb5383c897920aef31b42dd91da49be9",
      x"243cb5f543f6acba66104f3d87582fc4d8a67c555499159486a6dc00948daf9b",
      x"b843d402e1d618d038699aed15c39680e1c7f332597b75820c4eeeb5350aee3e",
      x"eec0531a10031f2d0ff6541bb34d1749ba0e373d11c5179368247f6af0b06b40",
      x"a006c7c11c91371e6080aa425ccea4ef5a66f4a36bf9a5600f36d4fd5c6d3d90",
      x"1bf5b6f90e1fba76d0a914c0ea4f6760a34953216bc39cc15d100aca7ea2682a",
      x"d1255678b649a89fb3f846514aaebb7211cf501f21e285a660e7779a52d4d566",
      x"0b8d3d1065180d4499b9a8c47057d715117fc196e813200e9b16004943b5ad36",
      x"5c7461001706a9573e3b07369c0c358d4f38583ce60caa83243556c950262cb1",
      x"1717d09db8a595b0b09af7c28bc6a3cf64731ba7d8363f00aa88d9851787ce33",
      x"2ebfe0b81e582af9ffda5bae0b119ee2f0ead7d209d4de1442c9c78ed666db5a",
      x"96ccbf8775211cfaa58e1444db9fce2102a72eaeee69cc99f1d5312b7d478ade",
      x"871e4dd055945902dfa180b20597d88956adff359f105b66bb4e6399ef567c88",
      x"f96a97a750cce3fd440ed33901be5ac632b686967de5a1767212cdec005f7bfd",
      x"306afed1e096f7b6b4201cf60295ba7f9492e67890fd425fe52e50d20caa2714",
      x"31f5ec03234adb88ee497b10acf242b335db6dc9cd1c9b91f6d2873dde9d8df8",
      x"4148afe3c3f50b4e5a23afa27e88070ff6dac6c91548614432ab658a41f3218b",
      x"6ae8e26abc160bc0b8c2c5cb1841ba5edf4678b25d72ba5d3e9015cb75dbbfd2",
      x"6e4e30d81fc0969916550d81dd3953f9b7ed177b7f5fb3fb25f8cf714dab07ac",
      x"dbd73b13bfda41ce35957e906899660b7e415f3a6ca023d9225047a02d539885",
      x"297368a199c836a28be13f17261e1b66b87db6545ea1e31c7efd7d9d989a3adf",
      x"5fa3619b4480c19499a52b85379dee418d5ce2439702099b09926ef3c3b17eda",
      x"5cb016b0acdffbc5eedb50076644842b43d819ea021cae280c28a1747294699e",
      x"f59940916594f8b443bbc0bfbb9898519199798721f2ced9fbf5364da1f660ff",
      x"406b26314fc972876def081781f5cb9447421c1a8a9c8c7b5268d2de9f408717",
      x"7de70eaebdb31bb00353cc00c4f2c84f5706ebece986db46bffc3b3f05ce7d33",
      x"29a0cfb8832e40ccdd4c8804e8711c0c3ca5af507e3e21cdbe10e4683cd94c56",
      x"6a75ea64df5f150956c883c446688fb28ca9f1a503bd7cd8db6b7cf21e4b8916",
      x"d0f65e85d98311cef3ddba8442acf16b9167189c9e012281963c8b53d4cf0df7",
      x"b7d76045984ebf006a42375b0bcf16e417f268a93f43ac56e62b8c258df3ecb7",
      x"9e50bab325e67f1518c16657e09e54f267d0259052846aa1548743c22f24ff5c",
      x"e6548544dab00ff4719d56b9ad7b93181a3eda25dbd6ff34369830623b1bacc9",
      x"584388b4bb7e2eb69cbd217999226e09252acd1f91624c73cdf8b26c2e8f0194",
      x"07b618c11478f1320ba5ffa59f8d073348b5794460bb5c3996ec304baf5fca80",
      x"74a1a25a6a03316f3410afc39f51272f81f2b1eac87816ae47482b4e83e139d9",
      x"2da98be76af58400997a6b6028124f488c54b2a727b4bb821e138750e0ae47ad",
      x"73a3ff75571beb3f24a7b4a5cbb8924a23fe12976c6e464dfe8c93bd462a070b",
      x"da6fe2ed3b3f6a85270f295b0e99b7f069e0a280d16aa1b8f2f01f0d7d0dc921",
      x"d1b984fe637ad7f5894f729293f23bcbf111de796da810235ae4aee684d7ffb1",
      x"7a8f25fe1dca259325d7e604d2386a2572b616c293fd239bf51c2a2c045d8d41",
      x"66fd924269dd8b3c0aa3efddd96f888919d7c7934c2b57a9418fa3e7a3dd9dce",
      x"f18156a3c7bd6a0284728dff48dccaf045e4941eac17672782a8af549bc3e116",
      x"f95af993ed8956e396a8242fa18755bde24babf43edac778e1a9e32be9712909",
      x"8b892f93ce1c98434585de5d0e77dc19aaaf8c0344982747cc76182a1fc25c7d",
      x"74ead417392af3cf0a7c88c29042a758545253a8ce3200923d62c4cf45355a62",
      x"866579052dc43bf276e40ceb5ca9da09fdf9d2a0cf7af7ee0f2262ca9cecacff",
      x"47ea07f4cb38df955095bab654f93f925b4c4f4588f06df0fe1ef5b8b3a8e547",
      x"e25078ef4ee6c16028bb2549745331ae44dbe9a98e441342022689d98a012f0b",
      x"4166786d2d73a641f43adf5379f1c8cdb3a2d6f92ffb2aca03ec78403065999e",
      x"e5d53fb9c85e151b06c5925c59616950d108f8a91483f9844a9f3c0ff7606fec",
      x"cf104fa3947544300839f0b3bf2b90ca3cf60e45d5bba60e3430c2107bebcbef",
      x"9a2100a81c88a867fd688d00a5623179e67ae600c78151114ba8b09d017c860d",
      x"0e39da9c5dd07ddefd05474244c28662a4183ec661ba13f1b91f0b4a543f9c25",
      x"03031bb1f7b550c048fc9ef48f0e01db2bc8eabd7ccc759928da52ca99d3479f",
      x"ed4c76346639fc030aee2e40867fcf5ed07418b357c97bf2cc499732dd573211",
      x"d4aab35b7b6b49c060a24f801e1b518044dbb125c07380367e3303405aa9884f",
      x"15d937da559fe67a77d7f32f36b6ef5ccb2ac880d104649c73ed701273c601fb",
      x"f6fd8a2483571741f9ab448401626052eead0da9efe21a66c58707edf2711b1d",
      x"282cabfd9ffc0428e639675dbd617afa01ea9a113c32c334e2745208088d2527",
      x"6f93332c73435b36b9b4df51b1e698e3b9be3f1bbe1e0323ef01ac4ecbcab99e",
      x"059014acba800bf67004a599b45667ad56e95c6f5b59562cc359c9911707a1a5",
      x"483b8d28271a59a075f8b50832d225aabd4dc0d517bb207dc7cdc6252da8d299",
      x"f32ef9156a68326445b798357476975c73340050d77baf9243581b2cbfa10a00",
      x"56bed234d49175e1e268c761470e1e0c1a05c382b5236f9f0fcd661900bcbe9f",
      x"d2a39cd7317043f9eafd597c00a2e0dd2f2f6709055e61aeffb4d64ee480f7f9",
      x"27995c8caabf732b266d13cc5a160bdfc29772f2432e20eb2291c60c8d2e31e5",
      x"dc704ff025ce34eeb2b399252b391bb16f367e791d410f5d996283b980519820",
      x"a07646af96b37b958a428ae684ee16b6db3f49cd94a39d7b1282dc6058e48643",
      x"221440e28cf07a16694248bec070c0e8a3807627c09d1d35fb5f5abc52cbdf0a",
      x"3e1ec0b8add19eb4263436601530783931806d834157a1b58a703047999f8c9a",
      x"ef41c2efb1387958ba70d7916b40a6950b12a9e7e9f98206e203f147866b38b1",
      x"002d9b3cb1ed63053288f523de643913b155565d391ca7799c5c1febe4380688",
      x"61c4d5b11ea8d903be8d5e9a12565ff9fe274d2b3a1c06cfdd43e5cba85f67ba",
      x"bf59fda3c8060754e126fb2bc846f63fc192a3e046f4db21f1dfb324c82aabbb",
      x"06bd628b431352533d8648606a49a27b7824b08cffdc97e13eecc0dce7455ae0",
      x"7b6511af5a1ad49b072d247457d48f70f0d24d6dbfa5fa5258aa4eb9bcc084fd",
      x"fc855f863c65d47ba54709f316023b2d2b7a38141ddb94060ec1db2e99a93d2d",
      x"972482bfcb35243738a155a2cc7c72ed6e43262e8dbd38e6afef390c98240819",
      x"6f17e207416ff42692ef72e538d1ec7187638fea6129e9f8b48ad99e7258acc4",
      x"9f1b2aefe36a16135f325d5a3441b45e229a4c3b692ebffe9e2f201970cf7ab9",
      x"4321366debcad798e43b1839ed822f117e6a7a0fb387e00845a0e6d6b5c1e220",
      x"0bc4b38632c0d93b3473764ffb505ab479d9e065f8a3728efc081943a4a629c4",
      x"2bb2bd4e9163613164a9a31b60fb07bf0b89629bc482c6c25f63e971af645b4c",
      x"106bb5a64a849adc9b059d06ce0357dffba4b0d6c4af370ad5b846cea4d07cf1",
      x"cdf1b9508023d15cb5c48518e1275996de735f9f9972a5493cd7fb172107d7d3",
      x"11a8fe9ca52ed6dd3ee6df4eb72b0595f836359d89705aaeb762113a4d121459",
      x"2336fff671454e9b9569ec30a03d076fff1790d97709ade57223cad7752abcd8",
      x"49b1f1cc99133395dcb53d057ef03cea32901eb29d60a27f7ee8cd861de305ae",
      x"879f8cbaf9518ba44230036925386111ba5ab091de73433cd22cf8f262b13e07",
      x"67f616737da3e728f58a2deb11f1d8562105a51da0ab3bdd9f3d3993b70d2816",
      x"002e79a47e02b5b146a1e0091adb491cf340fcb02333bc714bb39edd013f4e51",
      x"39e64a156121747a40d9bcf1b4c4cfef0aa019299dd2db1bc28ba4f73973e273",
      x"9cff86db1201db6e318eea3c2719aa90ab1dea81d01c3fee873c438d3ba4c47c"
  );

  constant RMATRIX : T_RMATRIX := (
    (
      "101001111001110111001110101100",
      "111000101001111111010110001111",
      "111011010001011100101011101101",
      "011000001100110011110100011111",
      "010111011111010001011000101001",
      "101100000010011010010111111111",
      "101010011100111101101100100001",
      "001101101010001110111010101111",
      "110011011010111111100011011101",
      "110010000110011001100011100010",
      "111000011111111001010101100100",
      "110101010011000101011110101000",
      "010000111010110101011101111001",
      "110001110110100110110001010100",
      "100100011111001001000111011110",
      "100001011100010001110011111110",
      "101011110010000110011001001110",
      "110111010011110100100000010101",
      "100001100000100011100000101111",
      "100001111000011111111010111110",
      "100000001101100101101010000100",
      "100100110001010011101010000101",
      "110101001000100001010111101011",
      "110001011110111111010101011001",
      "101010110001000101101100100110",
      "110010011110011011100010110101",
      "111111001101101011011001010001",
      "110011100011100111011000110111",
      "010001000000110010110011111011",
      "111011100110001001011111101110",
      "010010100101111111100010001001",
      "111110011011000110110100001110",
      "111001101010100010100010100010",
      "100000000011000011100000010111",
      "101101100011001110000101110001",
      "111111000010101111110011100110",
      "000011001100110011000010110001",
      "011101111011101111001011110001",
      "001010110111011111001111010000",
      "101100001001000001101101100110",
      "011011010000101010000110001110",
      "101100110110000101111101001000",
      "001001010111000111001111001010",
      "010010100011111111000011111010",
      "101000110110011010101110010101",
      "010010110101110000110000011000",
      "011000101110000111000110011011",
      "010101010101001010011111110111",
      "011111001100101100111010000010",
      "100111011111010010001001110001",
      "100001100100010001101100100101",
      "111111000110100111100111110001",
      "111101100101001011110101101011",
      "111110011110100100100001000101",
      "100100011110011011110011110000",
      "111101000101011001001100011101",
      "110010011110011011111001001010",
      "100001001101110001011101111111",
      "000100010010100000011011100111",
      "111100011010001110110110100011",
      "110100011010101111011100100001",
      "001100101100010000010011110101",
      "100010001000010110000011011010",
      "011100001010010010011111101111",
      "111000010000110100111101000000",
      "001110011000101010101101100011",
      "000001111000001100110000010010",
      "110101011110011001011010000111",
      "000011011010111011100110001110",
      "111010100111010110111101011111",
      "001110101011001101011101111111",
      "000110100111101111001001011100",
      "001000010010000110110100000010",
      "101100110100010011010101010010",
      "010111001000100000110100101101",
      "101100110001000010100010010110",
      "001100101000111111010111000101",
      "110011000000110011101000011101",
      "110010001110110001010010000100",
      "011100110001011100010001111010",
      "011001000111100101100010110110",
      "000000001100100110010010101100",
      "010011010110111000010010110110",
      "111011000000011111110000000101",
      "101100110101101001101111101001",
      "110111010011111100101000001011",
      "100111110111101010111000000000",
      "001001111111000110101100110011",
      "010111001000001101100100111100",
      "110000111001001010011011001001",
      "111100110001100111011100101011",
      "000011000010000111011001010111",
      "000110001110101100000011101000",
      "100001101011000001001011011101",
      "100000010001101001010110100101",
      "001000111001000110111001011111",
      "010111110000001001000100111100",
      "110010001000001010001110101011",
      "100000000110010101000011111110",
      "000111110110001011000101100101",
      "010010100111011111000011000100",
      "000100000011001001011001010001",
      "001011111101011100011100001100",
      "011111001001110000111101101011",
      "011001011000000111001001111110",
      "101111011101010011110011011011",
      "100011110010111110100101101100",
      "100100010001101101010011010111",
      "110010100000100000101010110000",
      "010101100101110000011000010101",
      "000100001011001010111111001010",
      "011001010111011010100100011100",
      "111111110011000000001011110011",
      "110010000011011010011011011001",
      "110010110100011110101100110010",
      "100010111000111111110110000000",
      "001101110001100000101111100000",
      "100000111111101110011100001110",
      "000110110010010101111101010001",
      "110010111100001101110000110010",
      "000110100000100110110001001100",
      "001010001000111100101010000101",
      "010011101010110001000100010100",
      "110110110011100010010001110000",
      "110111001110101000001010011011",
      "000011010001001000010101110110",
      "100100011000111001001101000010",
      "010110010101000101011111101001",
      "110111010010100110000111010011",
      "011010111001011110000000100001",
      "010001010110000101011000011010",
      "100000000110111010011011010001",
      "001100110001110110110001001000",
      "011100100000010110111110000011",
      "100010010110110100011101110011",
      "010000110011111010001110110001",
      "011100000001010011100110010011",
      "000010001111100001011111000010",
      "000011101011010011111010001010",
      "000010001100010101010100001100",
      "100110011010100011100110011101",
      "101000000100000100000001110110",
      "001111110101110000110010111000",
      "011101011010011100010101110100",
      "010011010111011111010101101111",
      "010001100110000000001101000000",
      "010010100011011101001100110000",
      "010111001101010010000011011010",
      "000110001011000110101111011010",
      "011110010101101000000010010100",
      "001001111011100101011001100010",
      "000101000101100011011111000010",
      "000100101101010110101101110101",
      "101001010010010110010100011100",
      "000010101001001110000110100001",
      "111100001000011010111111101111",
      "100001011110100110010000011001",
      "011110010000100100100000000111",
      "010111111000110111000001111001",
      "111000110000110110010110010010",
      "010101110110101001111111011001",
      "011011001111010100001010110011",
      "110000110001011110010011111111",
      "001101000110000110000110110011",
      "110111011011110100100000011000",
      "100100010011000110011000101010",
      "111111010101101000011011010110",
      "100100110101011100001100111010",
      "100010010110100110011001001010",
      "000111000010010101001110100101",
      "111000101101111100101000001100",
      "111000111110101000010101100110",
      "100001101010101001110010011001",
      "111010101011111111010001001011",
      "100100011011000010000000101010",
      "110110100010001100000101101000",
      "101010110100010001101100010011",
      "111000101011100110110101100101",
      "000001111111000110101111011011",
      "110110101100010100101000011011",
      "100100001010111010100110011110",
      "101110100011010001011000010011",
      "010011010100011010110100011001",
      "010001001110011000011110100011",
      "011110111001111100100001010101",
      "101111010000101010011000100101",
      "101101011001110001011010001001",
      "011100100011101010111001110110",
      "111110110000010101010010001001",
      "010010110001011110011101001111",
      "100110101001011101000001111010",
      "101001100010110001010000011100",
      "001101100011101111000001111111",
      "110111000111001111010001100111",
      "100000011101000101111101111110",
      "100001011101110110010100110001",
      "111110111101111000010101011101",
      "111011101100011011110100011110",
      "010111101000001100010101100011",
      "000110111000011010010101111110",
      "000100010011001110100011010010",
      "110100011010101111111001101110",
      "110111011100001000111101111111",
      "101000001100010001101010000101",
      "001001110110010000101010011111",
      "011110100000001100111010101010",
      "100011000111000000100011000101",
      "100011110001110111111001101001",
      "110111000010001101101001001000",
      "000100000010001001001100100100",
      "100110010100001110000111010000",
      "000011000000001011100100010011",
      "000111001001010100000011000000",
      "001101111110000011100111101010",
      "010010010000101100110000000010",
      "010111100011010110000111100000",
      "110101000100101010010101010100",
      "000001111111011010111100001100",
      "000111010111000110010000010000",
      "111100100011010111100000011101",
      "000101000000111001110101011111",
      "001111100010000101110101010010",
      "000000001000010111111111100011",
      "100000010111001111000011111000",
      "011100101100101001001110101101",
      "101111001100010110010110101000"
    ),
    (
      "111110101111001101100101110110",
      "111000101011001111011111011111",
      "100010100110101011110000000111",
      "000000000101011011010010111110",
      "110110100011010100011010110000",
      "100011100001010101001011111101",
      "010001111110011101010001110010",
      "000010110001011110111010101111",
      "101011110001010001010110101010",
      "111101010101101001101101000100",
      "000100011001011001011011010111",
      "111000100010111011001111100101",
      "011010100011001001011010010000",
      "111010000001011001110001100111",
      "101101011011010100001111011011",
      "111111101010000111110000101000",
      "101000100110100101001001011001",
      "010011100101011100111010000101",
      "100100000010000110011110011011",
      "101001010100001000111101100111",
      "010010001011111001100111100001",
      "010110111111000001001111000100",
      "100100101101111111111001101100",
      "011010110100011000001100101110",
      "111001010011110110001010000011",
      "001011100111110010011010001011",
      "110100011111110001001010101011",
      "111111010000101011110011110010",
      "100011011011000100001001101101",
      "110110111000100101000111111010",
      "101000000111111000001110111010",
      "100001001110110001100000101100",
      "010000011010011101111010110010",
      "111100000001001011111110111111",
      "110101011011101010111100001010",
      "000111010101001010111010010111",
      "011101110101011010100101000001",
      "111111000100011011110000010101",
      "010101001011010110100001010011",
      "101101001101110001110001110100",
      "010100011000101000111101111111",
      "001100110010001101101111011101",
      "000001111001000010100010000001",
      "010100000100000101111011111000",
      "100110100110100110011010101001",
      "010000000000001010001101100110",
      "011100001111001000101110110001",
      "110101001100010010010110010100",
      "101001000000000110000100100000",
      "101000011110110010111110100111",
      "111110100111011010000000001010",
      "110000110100100000010011011011",
      "001111010100111111010010101111",
      "110110001110110101110110110011",
      "111000110011101000010111000100",
      "010010000110101111111011010011",
      "111001010000011100111111010011",
      "000100011100011100111100011011",
      "110100010101010000110010010110",
      "111001011010100000010000011110",
      "111001001111101001101111111111",
      "110000100101110100100000010001",
      "111010011101000101000110000001",
      "111000100010101100011100000011",
      "111010011111100001001000011111",
      "111100111001110011101010111010",
      "111111100010000101101000111110",
      "010010101110011110011001111010",
      "111011101100101110111010110110",
      "010111110000110101111110111110",
      "000001011001010000010110100100",
      "100100101010101100000100110010",
      "101011111011110101110010111111",
      "100010101100001110111000100010",
      "000000010010000011101111000101",
      "110111011000001111101011001111",
      "010001010100010101011001100110",
      "000011100010110110000000110111",
      "000011100011001000000000111110",
      "111111000010110000110111110010",
      "001010011111110100110001001001",
      "000101110101001101010010101111",
      "000011110011010011000100110011",
      "110000000111110101110000101101",
      "011111001101101000011000001100",
      "000011001010111101110101101011",
      "011001011011100011010011111100",
      "000000110100111010100111111101",
      "111110000010111000010000111100",
      "100111011101000000110100101001",
      "001100111000001011011111001101",
      "001111010001101001010100100111",
      "110111011110010101010001101010",
      "101001001100101100011110011000",
      "100111111111110000010110111110",
      "101111011110010001001011100011",
      "101100111001101000111010100010",
      "110001110101001001011111010101",
      "111000111101100110101001101101",
      "110000101011011000100011011001",
      "011101001010010001001011001011",
      "001011110101010110110101001100",
      "010101111001011110011010111101",
      "010110111101001101001010010101",
      "110111001111011000110110111001",
      "100001101110101111101000110111",
      "011111111101010100100110011010",
      "000000000011001011110011101001",
      "001100101111011011000000110011",
      "111001000111000101011111111011",
      "110101110000011110000001111110",
      "011101111011100011010001010111",
      "010011101000011001111011011010",
      "001100111001010100001001101000",
      "011001101101001011100000001000",
      "011111011101101001010100100110",
      "100100000000010111111111001110",
      "010011110101000111011101110011",
      "011001000000111110010010000100",
      "111000111001101000101001111000",
      "010101111011010110000101010011",
      "010000101110010001101101001001",
      "100100100110110100101011110100",
      "110011101011111010000011101100",
      "110110101000001110101001111011",
      "100111110111110000111101100110",
      "011111100010001011000000110101",
      "100010011000001100101000000110",
      "111101010000111010001100100010",
      "001110101100111110110010000101",
      "110100010000100011101101010010",
      "011110111110001100111010101110",
      "101011101111011001110100000101",
      "110011111110110100110000011001",
      "001001011111000101101110100111",
      "001100000111010011100111000101",
      "110101100101110011011100001001",
      "010000100001000010010111011110",
      "011011111000010010111011101000",
      "101011010001101111101010111001",
      "110001000110100011110101100001",
      "100101111010010100111100011011",
      "010001010001001000100100000100",
      "011110111011111000110001110000",
      "111100001110011110011100011010",
      "100001000011111111101000011110",
      "110111001101101101110101000110",
      "010111111101111000110110110110",
      "011110101001110111100101101001",
      "001001110000000100000111101010",
      "000110101011010111000010100111",
      "010100100100110111100101100010",
      "100110011011011010010010110101",
      "011110001100101100111011101011",
      "001101111100000101100001110000",
      "100101110010100111011011100011",
      "001111100001001101101010100010",
      "111101110101101111010000101101",
      "001110011011010010010001010101",
      "101011011010011101010100101100",
      "001000001100101001100000100001",
      "011101000101110101010100011100",
      "001111111010111010011000010000",
      "110111100010011011010001010010",
      "101011101011000100000010010111",
      "011011001001101010111000110001",
      "001111010010101010100101011011",
      "101110101100001000010001111010",
      "011010001101100111011011100001",
      "110111001110001110000110110010",
      "010110000001100100101110110011",
      "000111110111011000000011101011",
      "110111011010011101101100111010",
      "110010010000011110000110010100",
      "011001010101100101000111010101",
      "100111110011111111010111011010",
      "010111000000110100100000000101",
      "001000100010001001000010111011",
      "100111100111111001011010100000",
      "011111101111100100010111011000",
      "110001011011010111001011001010",
      "010001101010100011101101101010",
      "010100011110111000011000100111",
      "011010011011110010101101001111",
      "111011100100011101111111100110",
      "111100101101010000101010011001",
      "000101101101110111001101001100",
      "101110101010010111100101100110",
      "100100110100001001111101100001",
      "110101111100110000001110010001",
      "011101100111010000110000101100",
      "011000010110110101001000100100",
      "011101010011110111101101101111",
      "101100110011010111101111100100",
      "011011010011110101000011001001",
      "100011010101011001000100111100",
      "110000011100100110011011101100",
      "110000000000111110001010101000",
      "111001110001000000000101100110",
      "101011011110001001100111001000",
      "001010011011100101010011000010",
      "100010000000000001101000011011",
      "111010011010001101111100101111",
      "101101101001001000010011010010",
      "101000001100010011001000000011",
      "001101110100110011111000101110",
      "110111011100000101001100100100",
      "001000010100111101000111111100",
      "010000111101100001000000111011",
      "000110110000000100111110110001",
      "100111000000010101000011011110",
      "010100000011011100001111111001",
      "110011110111111011100011110000",
      "100000010110110101110101101111",
      "011101110111011011000111001011",
      "001001000110011011011011001010",
      "000101001011000011110001000110",
      "000010111010001001110111100100",
      "100010111010100100011110000000",
      "101110100110110110110010011000",
      "000010101111001110101101101010",
      "000011010001011110010011110110",
      "000111011010100101101010011000",
      "110110110011110000101001101000",
      "100011111100000111000000001010",
      "110001101011111011110001100000"
    ),
    (
      "111001100000000011011101001011",
      "000111001001111011010000101111",
      "111100101011001011111111000111",
      "010001000100001000111100010111",
      "100101110000101001100001110110",
      "101010011001101010001011000011",
      "101000110110001110010101011100",
      "010011010101101110011101001101",
      "100101111101000101101111000000",
      "010011001111101011011010111101",
      "111011100011001100100100010001",
      "001101111101110111000101010000",
      "011011110010010001100001010100",
      "001000100011101001000110111001",
      "001100001001010111010000001000",
      "100001101010111001111111100010",
      "011011110001110000011010111000",
      "110111000010011011101110101101",
      "000000110110011110100110000111",
      "101000011010110011101100001110",
      "111100001000111011001001100101",
      "111010110110100111001101011100",
      "000010111101000100011101110000",
      "010110110111001101101000010011",
      "000101111000110000001000001101",
      "111101101011010100011111010100",
      "000110011111100101101111000110",
      "010010100100101011010001011100",
      "000010100101000011001100010000",
      "010000010101111010000001011011",
      "110001011011101111110101111111",
      "011000001111011101110001110010",
      "001000000101111111011010001001",
      "001001001110011100010110111000",
      "011011011010001111000100110111",
      "010011001110001010010000111000",
      "110000001100100110010101100011",
      "010100000100010100001101111001",
      "100010100111011101100001111010",
      "010001000101011000100110101110",
      "111000101010101100100101010101",
      "011010001111011000110110000100",
      "010101010000000101100101000001",
      "000110110110100011001011001011",
      "100111111011000011011110011111",
      "011010011010101101100111011110",
      "100011101100011001000101000100",
      "110010010011001110110000001110",
      "111010010011011001011110100100",
      "000011101101001100100001110001",
      "011010110111010110110011000100",
      "101001100001111001100011001100",
      "000100011001001001110011001010",
      "101000110001000100010000101111",
      "100000101011110100111111011100",
      "111001110111001111111111110010",
      "100111010011000000011001010110",
      "101010110011110110101101111101",
      "110111100101011000001100010110",
      "111000100100010000111111000100",
      "101010011101001110111101011100",
      "011000001000101001110011101001",
      "000111110101101011001001010100",
      "001101011011011110010110010101",
      "010110010110010000010000111010",
      "000000011001100100111110000010",
      "001110101001001001011110100110",
      "000010100100110011100110000010",
      "010001101111110010101011100011",
      "110011011111000110010011010101",
      "101111110001011000001010010000",
      "111111011100001101100101011010",
      "111101011111010011000110000000",
      "001101110011100010000100001001",
      "100110101101100001001111000101",
      "000010111011010000001011111001",
      "010000111101111100000001110110",
      "100100010000111100111101111110",
      "110110111000111001011101111100",
      "111100010111010110000010111000",
      "111001011100111110111011101101",
      "110110000111110100110111011000",
      "101010011010001000111101110000",
      "010100010101011011000101111110",
      "100100000000110001101110100110",
      "010110100110101011101010100111",
      "001010111100111001101011101100",
      "001011001101000100101111000010",
      "101010100001001101100110100100",
      "001100011110001100110111101111",
      "111111100100100011100111011111",
      "100000001100111101110010100001",
      "010100100000111111010100000100",
      "010101101110011011100011100101",
      "100011111001000100011100100100",
      "010111100010101111101000011001",
      "110111010110101100000111100010",
      "001011011001111100111100100010",
      "011101110010101101101110011001",
      "001100101110110010000100010111",
      "101101000111011101101000000010",
      "000100100011011001110010010111",
      "011010011000000000111010100010",
      "110110111011010101001110111011",
      "010100011000010000010010111100",
      "011100101010011010111000001011",
      "000111110111101100000010111110",
      "011101010110001110001010000100",
      "100001000101001100101001000000",
      "100000001110100010100000011001",
      "010011111111001110111110101001",
      "101100001110110011100010001001",
      "101011000000100101101100100001",
      "110010001100111010010011001001",
      "010111101001100100001000011001",
      "100101110110001010110100001000",
      "010100010001010101001011001100",
      "100100111001000001111001001001",
      "100011010011111100100000010010",
      "111000010101110100010110100101",
      "000010001010011110111000101101",
      "010011010100110010111110011111",
      "100001111101000110011101011001",
      "001010100100001101110100010000",
      "111101000000010000101001111000",
      "111111101101111101110011101100",
      "000110010010110010001101010001",
      "110101011011001001100011011111",
      "110001001110101101100010100000",
      "000101100100101000010001110001",
      "110000010110101001001010011001",
      "110110110000000101011011000001",
      "111110100111110111111010111011",
      "101010100011010010110000010111",
      "010001000100000101101100011110",
      "100110100011110011000010100010",
      "011000010001101010111110010000",
      "110000010111010000101101100011",
      "110010010110000011010110111101",
      "000011011000110111111000000110",
      "110000011110010100111011011000",
      "001011100000111100111111111100",
      "011010010010111010010010101111",
      "010011011000011011111101110001",
      "011011110101110111111001110111",
      "011111100101010110111111000000",
      "111010001000100011100101111011",
      "001010100101110110011100011111",
      "010000110101101011011110010111",
      "010011100100000011111101011001",
      "100100101101100011001111100101",
      "000011001110100011000110101100",
      "001100101100100011100001000001",
      "001110000101111000010000000001",
      "100010100100000100001110001011",
      "011010000111011000110100101011",
      "111101100101010100000001101100",
      "111110100001001110001000101001",
      "001001011100110100100010100000",
      "101001000110111001010010000011",
      "101001111010000101000111010101",
      "100000001011011110110000101100",
      "101110010000011100001011000010",
      "001101000111001011101100011101",
      "111110011010011110100101011000",
      "100000011010100011100001000110",
      "011111010010000111000000100111",
      "100000111100010000001100010000",
      "111001010100001111100110001111",
      "000011010101111100100011001100",
      "111010101001101100110100010111",
      "111100011001110101001010000111",
      "001101100111111100010010000111",
      "000110000110101111011100001100",
      "001011011001101011010110010010",
      "101101000001001001001001000110",
      "100101010101111100010101011011",
      "110101111100001010111111001001",
      "100111101110110110011101110111",
      "110011000110001001111111100110",
      "010010111101001110001000100110",
      "110111000101101111011000001011",
      "100110100010001000110000111111",
      "010001110001111101000000000110",
      "001110001101110101110010111101",
      "001101100110100101011101000001",
      "100100001001111000110000101001",
      "011101000101000000110110000101",
      "101010010000101000001000011110",
      "011100010011010110011110001011",
      "000101011010110101001101110001",
      "110111111111011000110101111101",
      "111111101010111011111101010011",
      "110111101111100101010000111100",
      "011101000010111000110100101100",
      "010000001111101011001101001010",
      "001000000010110010111100010000",
      "111110111011110111100101001001",
      "100101111111101100111011101100",
      "001000101010110110011011011011",
      "011111110001110100001110001010",
      "100000101001100111110010100101",
      "000001100010111010010010100101",
      "010110100100010001110111010010",
      "100101010010010000011001001000",
      "001011101010101001111001010000",
      "110101000010011100001101111101",
      "101001110110111110111010101101",
      "100001101010111010100100110011",
      "010011001101010111101011001101",
      "111000001010000010000010011010",
      "100001100010010011010101100100",
      "100110010010111011110010110110",
      "101100011100010100000101001001",
      "000110010001011001011011110010",
      "100111101100100000001110001100",
      "100000010011111011100000110111",
      "001101001010000001101110011101",
      "111011100000001000000001011010",
      "111101011000010100010011000011",
      "101010000110001000011110101000",
      "110011101000000100000001110101",
      "111100110111010011000110011001",
      "000001110100010001100011110000",
      "010011010010000110011001101000",
      "000010001001111100000001110000"
    ),
    (
      "001100110011101110111000110100",
      "001000110100000100010100010000",
      "010110110111111001100110111110",
      "110011100011000111001000101010",
      "111101010010000000111100010010",
      "100100010000101001011100010110",
      "101111000011111101100010101100",
      "001001000000001001110001110100",
      "000000100111011101100100011100",
      "101101000111111111010111001110",
      "111110100110100101000011001011",
      "010011000110101000100011000110",
      "000100000010001011001011111110",
      "001001001111000111100110101101",
      "101000011101101100100111000010",
      "001100101110000001011010101101",
      "111010010110101010111111010101",
      "101101010111101101100110101000",
      "101110001011011000001111011110",
      "000010000011011011000011000011",
      "000100010110110010111111001101",
      "011110001111000001000100100100",
      "000101101001001111011100111100",
      "010111111111101111001000000111",
      "101100001010110011111010000011",
      "010101110011010101110010100001",
      "101011001001001000001010101010",
      "101110011011110100101010110100",
      "011000000011011110011001000000",
      "100001110100101010100000101011",
      "001100010111101101001100000011",
      "101110100001100101101100101010",
      "111110000100010001111111110110",
      "001011100111001100001011101100",
      "010010001001101100001110100001",
      "001001011000101010111100100110",
      "100000001111111011001010000110",
      "101101110010000000111111110110",
      "110110111111100110010000100000",
      "101100010000001100000011111100",
      "000010101110000010111011000100",
      "101010101011001011010110111101",
      "011111010100001101101010100111",
      "001110101100110001101111010011",
      "010011010000001010100101110101",
      "011111100100001111011111111001",
      "000100100110101100101001100111",
      "110010110001010000101010110000",
      "001010000011110000010011000110",
      "010110101001001101110001100101",
      "000110110101011010011001101111",
      "011011010111101111100011111000",
      "100101110011100110010111010101",
      "110011000010010001111111001101",
      "111110001110010111110111001010",
      "100011100010100101001100011000",
      "001001001100001011001110001010",
      "110000111111001010100100100010",
      "010010110101101000111110101000",
      "111110111000000011001011000010",
      "010011010101101001001001110000",
      "101000111100001110011011110111",
      "111111110001111110111111010111",
      "000010001001100110000000001110",
      "101000111111111010111111110011",
      "011110111011001110010100011101",
      "111011010111111000101101110101",
      "101001101101001100010001001100",
      "110011100101100010110001111001",
      "001001000010000001101101100101",
      "101011100101101001111101111011",
      "111011100100000011010111101000",
      "100100011011010101100100010111",
      "001111011100101110101110001000",
      "100110101001100100100110000011",
      "011101100000100010010000000011",
      "110101110010000001001011110101",
      "111111110111101110101100111100",
      "011100000101110001101010110011",
      "011010010001110110000110100111",
      "111000000010101011001101001111",
      "111111001100101101010000001110",
      "001000100111101111100110010001",
      "100111000111111101010010110001",
      "110111101101110000001100101000",
      "101011000101111100110110010110",
      "110110110011110001111111100101",
      "001111000011001101100000011010",
      "010001101111100001100011101111",
      "010010110001000000110011111110",
      "111110000111110100100100100001",
      "110000011011111010100001101001",
      "100111111101000010101110010010",
      "101011000000011100011010011110",
      "011111110110001100010010100100",
      "011011001011101110011110111010",
      "010111101111110000110110100011",
      "100111000010010011100010110100",
      "100110011010011000101100101001",
      "111111110001001001101100010111",
      "010101100010111111011011001000",
      "011100101111000001000010000101",
      "011110111000001100000110110000",
      "110001101110001100100010010110",
      "010110011101010101000010011001",
      "101000100110000110101100001100",
      "110001100011010010110100010110",
      "001111011110011010101110101010",
      "011010110110100101100010010000",
      "100111010111100011001000001000",
      "000010101010110101110111111111",
      "111011011100000010101000111100",
      "111001101000100111001001011110",
      "110101000111000001010001001111",
      "111001100110101100111000110100",
      "111101011111110001001110111101",
      "101011010011100100110101110110",
      "100000000010010110010111101001",
      "111000010110100100101101101101",
      "001110101100110110101111011111",
      "011010100110111101001000101100",
      "001110100001011110101111000011",
      "111111011011000001111111011110",
      "111111010101111001001101111100",
      "101100000011110101111001110110",
      "011000010111111010001001110101",
      "011001110110000001000101101010",
      "001010000010110000100001110011",
      "100100000011100101110110101110",
      "110011010111101111110100101000",
      "110110110101000100010001111001",
      "100001110110111111011101100111",
      "111011110011100100110010111001",
      "011100101100101011100111011010",
      "101111101001010100101101100011",
      "101101111100101011001000000100",
      "100100111011011000001100101000",
      "001100110011010011001111011001",
      "100101110011011010010011110101",
      "000001111010101110010010101111",
      "111101101011100001110000000001",
      "001000111110100010111111011011",
      "100011100101111010110010111100",
      "010011010010111001111100000100",
      "011010011000001010101010111111",
      "100110110111100110101011001000",
      "110011110010111111111010101000",
      "111010101110000011011110111100",
      "000001110100011101001101111110",
      "100101101101110101101000001010",
      "101001100000011000000010010101",
      "010000110101011110001010111110",
      "110001100110111110000100011101",
      "000110000001011101100100111110",
      "101100111100000101011111011101",
      "101101000010001111101010110111",
      "101111001011111000000001110111",
      "000111100010010111000101100111",
      "100011001100000011000010011011",
      "000001100101111011101001111100",
      "010001100111110000011101110000",
      "101000010100000011110000110010",
      "101100100010001010000000010000",
      "011001011101001111110000101001",
      "111110001110011011011001101001",
      "111101000011010011010111110101",
      "110101101001010000110101011011",
      "101100110011111011101001011000",
      "101110110110100001110110011100",
      "111110110010111110100101100110",
      "100111000110111011011000100011",
      "110101010111000111010101000110",
      "110110000010101000011111111000",
      "001111001100010010111000110110",
      "010010001001111111001010111100",
      "110000010011011101101001000101",
      "010101101110101100110100010011",
      "011001111111100010111100000001",
      "010110101000110100011100101011",
      "000110011001100000001100000000",
      "100011011011111111001110100000",
      "110111001001101011011111001011",
      "110101010111010001000110011010",
      "000010001011001000111010000001",
      "100100100011110111000011111010",
      "101100001100101010001101101110",
      "001011011011110100101110111110",
      "111010100001110100101001010010",
      "111110110111001001010110010010",
      "011101110101001111001101111011",
      "001010100011101101101000011110",
      "100110110110101100111111001110",
      "000001100011101001011110100011",
      "110100011001010111101011000001",
      "011001011111101111110000000111",
      "100001001111110010100001101111",
      "010110111110111101001101010111",
      "000010101101010110110110111000",
      "101100101010100010010011010101",
      "111101111001100101101101001011",
      "011111100110001110110100010010",
      "111011101000111101011110000100",
      "011010110000110110110111111000",
      "101100100101000010101001101110",
      "100110010110111111100010000111",
      "111001101110101011111001011000",
      "001100100100101111101111110000",
      "000100010100001010111011010001",
      "001001010111000111001111011000",
      "111011100110100101011001101000",
      "101011000001111001111010010000",
      "001110000101111100010010111100",
      "111100001010100100000010111001",
      "101100111011011100101100111110",
      "010010110010011110000001011010",
      "101101110011010101100011011011",
      "101001101001100110011111011110",
      "000010000001101010111001001100",
      "010000111110110101101100111100",
      "101001101001111111111001111000",
      "000110101101010010011110001110",
      "101111100001110111101011101000",
      "101001000011101001100011001111",
      "001110111100111111001010011001",
      "101110101100011011101011101001",
      "011100000010010001011001000000"
    ),
    (
      "011100001000110111110001010010",
      "100010010001000100100000011000",
      "000011100000000000001000110010",
      "000010001000110111100100011010",
      "101010101000011000101110001011",
      "101000101011111100011001011111",
      "100100111000000110100001111111",
      "110100010001000011110011000100",
      "000010101110100101100010000001",
      "100000000011100101111111111001",
      "110100000001101110101111110101",
      "100101011101001010011110010111",
      "110010101101001101111101110111",
      "000111101111010000001101101000",
      "000010000111010001101010110011",
      "100011111010000111011011010111",
      "100110001011000110110110000000",
      "011110010100000111010110011000",
      "101101110101101110011110101001",
      "101010000000110111000010010010",
      "001111110100101010010100000101",
      "000111110011100011110101110001",
      "010011110011101110010011111000",
      "001011000100100100100001001110",
      "111000100010000110100100000101",
      "111101110010011011001100010010",
      "101110111000010100111000010011",
      "111111000100100000011110001010",
      "000110001111101001101001100101",
      "110111110101110011011001111000",
      "000001001010110101001011011101",
      "101010110100001111100110011000",
      "000101110000101001101110011111",
      "010000000100111100101110111101",
      "110010101001010000110001000110",
      "010111000011000011000111001011",
      "111100010100101100101001101101",
      "101101001010000001001011110001",
      "100101100011111000001001111010",
      "000000011001100101010011101110",
      "110010011000001101101000010001",
      "110100000000111101010000000010",
      "110000110110000010100111011100",
      "011100010001111010100011100101",
      "101011010111110000110011011001",
      "101110011100001010000001010110",
      "101000000100101011101001001101",
      "000110100000110000010000101111",
      "100100011010110001100000110101",
      "001100011111101101011111111001",
      "111001001110011100110001101111",
      "111010011011011111001010100011",
      "100001001110000001110001101111",
      "100100010010101100001001010101",
      "011110110100010100101000111010",
      "100110100111101101001011111011",
      "101100110011110001010100010000",
      "101110110111100010110111110000",
      "010111111010011001101011110000",
      "100000101111011110010001000001",
      "111011001001001000110001100110",
      "001001000100100101011101010000",
      "110011000001100010000001111001",
      "001110101111011010010001100100",
      "001011111000111010011110110111",
      "000110100010000100101001110000",
      "110011100000010010101011010011",
      "100111001010001010011111000101",
      "010111010101110000011000011110",
      "000111101001101010110001000011",
      "110001100110001000111110100110",
      "001000000010110010101001011100",
      "000001010010000110111101100111",
      "000101110000100101110011011011",
      "110001010011111000000110011000",
      "000000111101100100101001010000",
      "001001011100111100001111011111",
      "000001001001111110001110000101",
      "111001111000001101001010111110",
      "101001100101101010101110000000",
      "010100010011100100101111111110",
      "001111010111010100110010101101",
      "100111010001011010000111100110",
      "111101001100111101100111011010",
      "000010010000000001101001010111",
      "101110001011001011001001010001",
      "010000000101111010111000100001",
      "000011111011101100100111001000",
      "010111011010011011110110010100",
      "010000111011001001110000101101",
      "100100011001111001101100110111",
      "101000000101101000100110111011",
      "111011110111111110100000110001",
      "000101000000101000110111011110",
      "110010100011001001111011000101",
      "001010111000001100110100110010",
      "100001001110011100101101000010",
      "100111010110001100011000100100",
      "001000110101000001011011100111",
      "100001001101101000010111100010",
      "011011111100010010011011011011",
      "001011010101101001011101111010",
      "000100100111000111000001000011",
      "101110011001110100010000000101",
      "010010110101110101111110101000",
      "011100001001110110111001011011",
      "100001001100110101110011100000",
      "000111110011001001011111111010",
      "011001111110010111011000001101",
      "111010000010100101111100101101",
      "001010010010110110010110000100",
      "101010000000111001101110111011",
      "010110011011011100101001000010",
      "111100000110101111001011010000",
      "100101100101111100011110100001",
      "010001010101101010101000100110",
      "111111001000110000001111000000",
      "110010001001001110101111001101",
      "000001000011110001101001100010",
      "110000001011110111001111011001",
      "001001101100110000010011001111",
      "011000001011010011100100001010",
      "110100110000111100011001010101",
      "000001011101110000010111101011",
      "101010000110100000010010001110",
      "101000010001101100010101011001",
      "010011010101011111000001010100",
      "000001110111101010001001101110",
      "101001111000010110011101111101",
      "001011010101111001001101110101",
      "111010011100001101011011110000",
      "001101100111000000011010011111",
      "101101010010101111110011011101",
      "111110100011000010001100110101",
      "010111010010100001001000001010",
      "011011011001110010111111000100",
      "010001000010000010100001101100",
      "100001010011111111010001011101",
      "000011101111011001001101000111",
      "111110111011111001100010000100",
      "110110010000001110101110000010",
      "000000110000000000011001111010",
      "000110101011011000011000000011",
      "010000111011101001010110000000",
      "001010110101110101101001011100",
      "001110111001000111110001000100",
      "111010010010010110010000010001",
      "010000100001011000110110101110",
      "111000110100010111011011110010",
      "101100000111011100111000100010",
      "111111010100110101101010011000",
      "100001101001100000010011100000",
      "011000111011011011101000010000",
      "101010110111000100011010100000",
      "011100110100110101001001010000",
      "011000101110111100010010110000",
      "001101110010010000101010110100",
      "110110110101100100100001101011",
      "100010000111110111010011110110",
      "001110010111110010100111000011",
      "000011000100100100011100000000",
      "000000101100001000001001100011",
      "001111011110110100001001000100",
      "000101001101111001111110010000",
      "011011000011110010101000101101",
      "110101000011101111101111010110",
      "100011010000000010111100100100",
      "001101110011110101011111000100",
      "110000100011001001101001000100",
      "000001111111111010111110100011",
      "100000000000011101001101001001",
      "110101011001000101001001010111",
      "000011000001000100011011000010",
      "101001100101100001011000101000",
      "001011010111000011000100001011",
      "001100100101011111100100001000",
      "000000011011101000101100100111",
      "001100000011001100100000010010",
      "110000001010111111100111010010",
      "010110110101110111010010010000",
      "011010101011100110101001101011",
      "100111100110100010001011011111",
      "011001000110110101100011000010",
      "100000110101001000001011111011",
      "110111101110111011010001000001",
      "100010010001100101010010010111",
      "001100001001001110001100011110",
      "111100101110011101011011001110",
      "110110011000110011111010010010",
      "000010111000011110101011100000",
      "010111110101100011111011110000",
      "011001010111001111100011101101",
      "010111010011101101111111010101",
      "000111110001111000110110001011",
      "101100001110100110010010011010",
      "101100111011100000011011011011",
      "110100110011100011111101001010",
      "010100101110010000000110000110",
      "010111100110001000100010100111",
      "001001001001001111101111111110",
      "001100011001110000010101111111",
      "110110011101110001010001011000",
      "111000010001010101100101010111",
      "111111011011001001010011010010",
      "000100111010000100111011001110",
      "111111001010011011000010000100",
      "000111111100101000001100010101",
      "001101111111001001101000001100",
      "000100000100011111001110010000",
      "101110110101110010000010111110",
      "100010011011011011011000110100",
      "000101010010111100010100110101",
      "100111100111101000101100010110",
      "010000111000111101011101000100",
      "000101110001010000000011101010",
      "011111111000100110101111011101",
      "111000100100111100000001010101",
      "110000100100000110001110100110",
      "000110101001001010001000010001",
      "110111011011111001011101010010",
      "110110110111111111100101100010",
      "100111010111100100010010101111",
      "101011111101010100000110010110",
      "000110110101101011011000111100",
      "100000000111100101001010100011",
      "111110101110111110001001000011"
    ),
    (
      "110101001001010100111100101100",
      "010011111101000100111111010100",
      "100100011011101011001010010011",
      "000110000110110011110100001010",
      "100011101000001000100010010011",
      "110001100100011011100001100001",
      "100000000110110010011010101011",
      "101100001100110011110100010001",
      "101100010001101010110100010110",
      "000001011101011100011010100111",
      "010001011100111010100101011110",
      "010011110010111010010010010011",
      "001100110100111010101011001011",
      "100110011110100011110101110111",
      "011010110110000100001000001010",
      "111100111000011111011101110001",
      "101000001011111001111100100000",
      "010111001000100111111000010000",
      "001010000101001110001100110010",
      "100000010111001101110001100101",
      "010011110001110111011001100110",
      "100010000101000101110101011100",
      "101000110000111010101101010000",
      "011010000010011110001111010011",
      "101011101101001101101011000010",
      "111111001010101110101001010100",
      "001110010001110011110010010110",
      "000100000110111100010110000010",
      "111111111101111000001110001110",
      "011110101101101000110111111011",
      "010100101100101100110000110110",
      "000111010111010111101011001111",
      "011010010000111011101100010001",
      "000001010111010100111111010111",
      "111010101011100001011101110100",
      "101110001001111101011000100001",
      "000110010000101011010001000010",
      "110100101100000000001010010000",
      "000111101001001110110111100000",
      "111110100000110111110101010011",
      "101000110111100110101000001000",
      "101110111111001111000001100100",
      "000110011110001110100100010110",
      "000000010001000011011101100110",
      "110100101111101101000100100111",
      "001001001111000000000011010011",
      "001000000000110011100111001100",
      "001010011001100001101111110011",
      "000101001010001011100000100100",
      "101000001001000000010001110011",
      "000110011100111010010001100100",
      "001111011110010001000011001111",
      "010100011110110000111010001111",
      "111101100110101100010011100011",
      "101100000000101001111000101001",
      "010001001000111010111100011101",
      "101000101010110000110000011000",
      "010001100010000011101101111111",
      "111111101110111111111001111100",
      "111100111001001000100110110011",
      "010111011101110111001000010010",
      "010110001000110111111110000000",
      "001111101000000110111101111100",
      "100010011101011010110110010001",
      "100111001000001100000001011100",
      "111000111000111101000110100010",
      "111100110110101101001100111100",
      "101111001101100010000001111011",
      "100111100101011111101100100000",
      "100101011101011011010100011111",
      "110000011010101001110010100111",
      "100010010010000111001011011111",
      "110000101111010010001111100101",
      "011000000000111010010010011011",
      "100010111010101000111110011000",
      "111101101101111100001100000110",
      "110110110000110001000000000001",
      "110010101110010001011010001010",
      "111000010001100011001000000100",
      "110101001110101101011111001001",
      "010000100001010001111100001001",
      "001000000111101011000101010000",
      "001011000010011001010000011101",
      "110000001001111011001100011010",
      "111001110101000011001101001110",
      "110000011011000100011111000101",
      "011111111110101111000010001101",
      "111001011101100111000011011001",
      "100000111111001110111001100001",
      "001010010111011000110100010110",
      "011001010000000101011010100000",
      "111111000111010101111010000001",
      "111111110101001101010001010000",
      "011001111010010010100000100100",
      "110111000000101001100000110010",
      "101000000011001010100011110101",
      "011101111110010110010110100001",
      "100011101011101001010011010100",
      "110001111001001111010011101010",
      "010010100001111001001001101110",
      "010100010100011010000011110101",
      "111001100101010111000101000011",
      "010111000110101001000101100100",
      "000111011000011110000001100011",
      "011000111010001111000100111100",
      "001110000010010010100001010001",
      "000001111110000110111110101111",
      "100100010101001101001011111100",
      "010110001000000100011011001001",
      "001100100001111101110001000001",
      "011001011101111101001001111011",
      "100011000011110001010000100000",
      "111001010000000010000101100010",
      "000110100010110010001100111010",
      "111101110001111110101011110100",
      "011001111000000011001001011000",
      "010101101000111011010111011000",
      "100100100000100001100001101110",
      "100000010111011001011011010000",
      "001011100000111010100011001100",
      "101010001001011100001110111100",
      "000011100010111111110110000011",
      "011000101101110000111000101110",
      "101100001100111100101001010111",
      "101101001110010101000011101010",
      "001010000110010000111000000011",
      "101011110011101011101001011011",
      "100111101000111011101000110001",
      "011101111101100101101010111110",
      "001111001111010010010011000010",
      "110100001011111110010000111101",
      "111110100111100001010001111101",
      "011100000001101001010010001111",
      "111111111100101000010111101010",
      "001001001100111001110110111101",
      "101010110000100000100111000110",
      "010111111011011011011011001000",
      "111010001000111010100011010101",
      "101000011111010101110000010100",
      "010110111101010011001111011100",
      "101100111001101111111110101011",
      "000111111000011010110110000001",
      "010110010001001100001011000110",
      "110110010100010111100010001001",
      "100111100011101010000000110000",
      "001011111011000101101011111100",
      "101010010011000011101111110110",
      "011010100111101000001100000011",
      "110011001111001100101001100111",
      "100101010111100110100010100010",
      "010010101101000101000110010011",
      "010011010000011110000000101111",
      "101110101011100100000110000011",
      "111100001100101001011000111111",
      "100000110011110110000011100000",
      "010010011101010101110110000010",
      "101110110001001011100100101011",
      "101010011110100110110111001000",
      "000101110011011110110100101111",
      "010011111110100010011011000101",
      "100100110100001100101000000110",
      "101111110100100100101110011001",
      "101100110011110101111011001111",
      "101101100100100100011111101110",
      "101111001101111111010011011010",
      "011111100010010010101001100000",
      "111100011100110010000100010100",
      "101001101010101110010011010100",
      "101000100010001011011111100101",
      "110101100101000100110001011110",
      "111110001111011010110110111011",
      "101110100101000001000101000001",
      "110100010001000000110111011010",
      "101001110100000001011110110101",
      "100100011001101001010111110011",
      "100101110000110010000001011011",
      "010101111011001011110001011010",
      "101111000011110101001011101001",
      "100000010010001101111001011100",
      "001100001010001011111100100100",
      "000010100010111010000100110010",
      "110001011110111101100000000101",
      "011100011111001101001110010111",
      "011000100101100100101110000101",
      "011000011011010111101111000000",
      "110001101001010110011110101001",
      "111101100001101111001010111010",
      "110110101011011001000000110011",
      "110101001111101111011100110100",
      "111101101001100111001110100101",
      "001011010000011010001111110010",
      "001010001100100100101010011001",
      "100000001011010100000011100110",
      "101010110010001010101110011110",
      "001011111001001000101001000111",
      "110110110101111101101000010000",
      "011101011110011110111011011010",
      "001101110010000000110001100111",
      "111110001011111010000111001001",
      "000100111000110000111111101011",
      "001000010011011010000100010000",
      "000010111100010001101000101010",
      "110110111111100100010001011101",
      "110011011111111010110011111001",
      "111010101111111100000100111100",
      "001100011100111001011000101101",
      "010110011001111111001000000111",
      "100101000111101010101000101010",
      "010100011000010001000110001100",
      "111001000001101011101110100001",
      "101010010101011111010100011111",
      "000100110010011111100010100101",
      "110101110001101000100011011101",
      "101101000001000101011011010000",
      "101010011110110000100010000100",
      "111101000010111010000101001110",
      "000000100010000100111100000001",
      "110111110010000100001010001111",
      "001111001001000011101100000011",
      "100010110111110001001001001110",
      "000001101101100110000010111000",
      "001101111001011011010101111010",
      "111011111111100111010111101011",
      "110011111010110010100111100000",
      "101000010001111011000100101100",
      "100111100111001100011101110000"
    ),
    (
      "110011000101010111001111010101",
      "111000111010110110001101100111",
      "110010001000110001100001010110",
      "111110001110001011101011011000",
      "101110110100011000111110001100",
      "101111011011101100001110111000",
      "100000010000001100100100110001",
      "001110011010111010000101111110",
      "001010100000110101010111101001",
      "100001000101101010010101011001",
      "011000011111111101100011001011",
      "011110110100001110101101010011",
      "010110000101010101001111001100",
      "010111001101111001000111001000",
      "100101000000000110000101101101",
      "110000110000101101010010010111",
      "101000111101110010100000101011",
      "010101101010101110001010110100",
      "101101010111101010011101111101",
      "000110101010000110000101011110",
      "000100000010100110010110011101",
      "001100010001011110101101011001",
      "001010110111010111010001110101",
      "101011110101110111111011000100",
      "110100011111110101011110001011",
      "100010000101010101000001100011",
      "000001010010111000100001001010",
      "110110001011010100010010111100",
      "011010000111011111001100000100",
      "001000001000001010101110010010",
      "001111010001101011111110000011",
      "011111001010110100111000100011",
      "000000111001000001101111001001",
      "111101101100101011101110001101",
      "110010100101011000000110110110",
      "000111111010101110100010111111",
      "011000011010101001000110001011",
      "001100011001100001010000110111",
      "000111000101110110111100001111",
      "000101101101011000000000110011",
      "001000001101000100111011000000",
      "000011110110110111111110110001",
      "111101001001000100111110010111",
      "111000110111111010111111000111",
      "000001001011011011100100101010",
      "100011011000111100111111001011",
      "011010101000010110000100111011",
      "101000101011011110101100101111",
      "001010100101100101100001100001",
      "001010100000010001010010111001",
      "011111010000010000001000110101",
      "111111110011100001100101010101",
      "101000100011000010001110101111",
      "101010110011000110001001011011",
      "111010011000100010000111001100",
      "111110000011111100000110100001",
      "100010101110001010110100010110",
      "001011000101100111100000111011",
      "101101110110011101001100111011",
      "111001100011101100001010110100",
      "100110001101011001010000001011",
      "110000011001101111110010001111",
      "101100001111010100110011111100",
      "001011100100000001100100100100",
      "001100011110100001010101000110",
      "100101010100100110100110011100",
      "100000111001001110010010001010",
      "000100001001001010100100111101",
      "110100100000100011100111010100",
      "010001010100100101001000100001",
      "001111001111101000110100101011",
      "000110010001000010001110000100",
      "100011010101101100100101110011",
      "011000011010100001010000001001",
      "001000111000011111010100011101",
      "010100111011100111100110010111",
      "111101110010110101110010001010",
      "011000011001000110011001100001",
      "010011001101101011011001100000",
      "100000000011111000100101001101",
      "010101110000010001010100101010",
      "000010010111001110111111001110",
      "000010110111001110101001101100",
      "100100001101000001100110101010",
      "110101001011000001110111100100",
      "100011101101101011110110100100",
      "100000011011111101001101111001",
      "110100000000110101100011100011",
      "111100110111111101101100100111",
      "010011000011111110001001010010",
      "101010101100010000110111100101",
      "000000101010111010100011000000",
      "011110110001100010111110110111",
      "111110100110010110011001110000",
      "101101001110011010000110111111",
      "010000111111111110110110010010",
      "000000011010110010011011001100",
      "111110110111100100100111000000",
      "111101100100101010000100111001",
      "101000101110101101011110100110",
      "001001011100100010101010101011",
      "110100010000000110001111010110",
      "101100001101101101100010110101",
      "000101111010111001011101011101",
      "000001100110010101001110111100",
      "001101010111001110111001111010",
      "111100101010101010011111010000",
      "000010110100111100111001100001",
      "101110000010110001001100000000",
      "100011010100011001010011000010",
      "110001110011100001000011010111",
      "011110110100111010001001011111",
      "000111011110010011100110101010",
      "101001001010001011101001110111",
      "000010001110100111111111100101",
      "001011101001001110110000000111",
      "101110001111111011110001111101",
      "001100110010110100000000100111",
      "110101001100000000110010110110",
      "011111111011101011000000010110",
      "101110000010011110011101100011",
      "011000100000111011011110000000",
      "010001111000000100101100010000",
      "110100011010101111011110001011",
      "110000001001110100011101110010",
      "101100111111010110010111011100",
      "111011010100100010111010101111",
      "110011111111111000100110111011",
      "111011100100100001110101111100",
      "010001001100110010010010100101",
      "110000001111001101001000100010",
      "110101000110011100001111100000",
      "010001001000111000100110110101",
      "101010010110011000010001100010",
      "101000001100111001011101101000",
      "011101110100011111100100111100",
      "001110101101110101001010000101",
      "101111001011011110011100100110",
      "010001001101010010101000010111",
      "001001101100100110001101111001",
      "111110001011110001010110110001",
      "000111010111011010000000101011",
      "011001001011011011111111001101",
      "101100110000101011000101111111",
      "101001100100100111100110000000",
      "010000010001100110101001010001",
      "100110100100111100101101011011",
      "010001100110011001100011011001",
      "001011100101011100010110110111",
      "010011101100001111110111110000",
      "110000000100010111001001000001",
      "010110101010100001110000100110",
      "000000110001010001100101110111",
      "111111111101101101100110000001",
      "000010000111010000110001000010",
      "110101111000110111100111111010",
      "011100011101110001110011000000",
      "101100101001101110000111000000",
      "011111011011110100101010001010",
      "110010001001000100000001000011",
      "100110100001101001111110011111",
      "001111011011000001101111111111",
      "001000100111000100101110011110",
      "100111011000100110101100110010",
      "011110011001000010111001100100",
      "100011101000111010110011011010",
      "010100001010010101001110011001",
      "010011001101000111010110011010",
      "111011000011110000110010010100",
      "011011111000110000100011010011",
      "110011110000110100111101111010",
      "010100111001110110000001010000",
      "110100110100010100000010110001",
      "100001111011000011111111100110",
      "001111000101000011011111100101",
      "111001010010001101110011010100",
      "010011011110011010001000001001",
      "001100010111111110101101100001",
      "111001000001011011101010100111",
      "010001101000001000000011011100",
      "101011101010110111011000010111",
      "001000001010000000011110110111",
      "110011011010101101000110001001",
      "011110001111010101011100111110",
      "000100000110011110101001001100",
      "011110111110100010100010110001",
      "101111110001100010101000011101",
      "101011001001100010000110010110",
      "111100110011011100101001011001",
      "000000000100101011010010100011",
      "011110100101111111111011010111",
      "010011101011101101101000001011",
      "100010110000100110000000100001",
      "010011010110010001100100100101",
      "110110000000101111000001111110",
      "001001011010110001011011001011",
      "001101111110101000000100110111",
      "011011010011000000011011101111",
      "110101110010100101100111111000",
      "100011101100101000100100110000",
      "010100101011010000101100011111",
      "111111010111001111100110011001",
      "000010010011011100011100111100",
      "001000100101110101001101010000",
      "111001110011100101100011000001",
      "100001111011101000000001010101",
      "001111111100000000111001011001",
      "001001101011000010100111000011",
      "010100011010110000111011010101",
      "000000111100110010110110010001",
      "101001011000110001100010100001",
      "010001101101100100010001000101",
      "101000111010000111011000000101",
      "100010001010000000111000001001",
      "110001111000011110101001101001",
      "110011111111011111011110010100",
      "001011101111100101011001111010",
      "100110011101101010011000101110",
      "000111111011111001100001000011",
      "101000101110100010000000101000",
      "000110001011100100110100111010",
      "111111001100011011111100100110",
      "100111000100111111101001000010",
      "010001110011101111101000101100",
      "000100101101101010111110110010",
      "000100000010111010101111100100"
    ),
    (
      "001001101100110000011100000101",
      "101110000101001000000011111111",
      "001100100011000001100000000111",
      "010010000101011000101100001000",
      "110000000000100111001011010001",
      "001001001100100100001110010010",
      "101111110110010011011000111100",
      "011010010101000001111001100000",
      "111011100101111000100100100000",
      "111011111110001101111110010111",
      "101110010010011111101100100110",
      "110110110101101010111101110000",
      "110111000101111111000010110100",
      "011101010100110011110010101011",
      "000111101010101110101000011110",
      "011011100001100100110001100111",
      "001011101100001001111110011110",
      "011111010001001010011101000100",
      "011110100010101111111011000011",
      "011100110001110100101011101000",
      "110000001101011110110111010010",
      "110010010110011101010110010110",
      "001001000011001010101110111111",
      "101000110110001101001011001011",
      "000111101000000001111001100010",
      "111110001011110000010011011001",
      "100010001010111011001111001111",
      "000011110011111111000111000110",
      "100000001001110000000111100111",
      "110000011101101100001001101000",
      "011010011000101011000010011111",
      "111110001101000100000010001111",
      "110001110111001011101001000100",
      "101110010100001011010100000000",
      "100110011110000011111011010100",
      "001011010011010110010011011110",
      "011011100001010000000101101010",
      "110010010010000100011000011000",
      "100000011010110101011110000100",
      "100100001011011101111111100111",
      "110001110001000010100001001001",
      "111011011110100111001001011110",
      "101100011110011011101110101101",
      "110001001110001001100010110000",
      "010011111011110100100011011100",
      "001111000101011100011001001011",
      "001011000101001101100100000011",
      "001001000001101001000000001111",
      "000101010010001001000011110011",
      "111001001110010110010001111001",
      "011101011001101010000000010011",
      "101100101000010111110010000010",
      "101110000001110000111101111111",
      "101101100010011100100011010110",
      "001011001000110100000011010001",
      "010010010101001110000010011100",
      "101000110111001110111111111000",
      "101100011011000001000010010011",
      "110000001101110100000001000010",
      "010111011011100000011000010001",
      "011011100001011011011001111110",
      "000000100011111110111111101001",
      "001001000011111111101100011100",
      "001110001110101011110110000100",
      "110000100101111001101100111110",
      "111000101111000001010001000010",
      "110011001100001110000111000001",
      "110100011011001110011111000100",
      "010010000001100100000101000011",
      "000101101001000111010000011111",
      "001010101100010011111011110000",
      "110011011000101010010011000101",
      "000000010110000010110101000101",
      "001011001110000011001001011110",
      "000100010100110010010110100110",
      "001010110111101000100011111000",
      "100001001011110111000000011111",
      "101000110011001110001000101000",
      "001111100010111111010100111010",
      "110011101110111000110110111011",
      "110100101011101101100110001010",
      "011101010101011111100110101001",
      "000110101001110101100010010001",
      "100011010101111111011011110110",
      "010100011100010110101100011110",
      "110001101101000001011000000110",
      "010010110100010110110000001000",
      "111010111001010110011011110010",
      "010000101110010001011111110101",
      "011000011111011110001011000110",
      "000110010001100101111011100000",
      "101010010001000011111000000011",
      "111100010000011111001101000001",
      "011000011010000010101000010110",
      "000001011110110101001110101001",
      "001000011110110010101010000110",
      "001110001011100000111011001100",
      "011101011100011110000101010110",
      "000010011010111010101111011001",
      "001000100001011001111101111001",
      "101000001100011111100111101100",
      "101001110011111001101000001111",
      "100101110101111101101001110000",
      "001001011000101110010000100110",
      "100111000000000011000010001111",
      "110100100110111000011101000000",
      "011010101110110111000110110111",
      "101101001011000010010101101100",
      "010110100000010101011000111111",
      "111100111100011001001010111101",
      "111011101100010011111110000001",
      "100000100010001100110101000010",
      "001000011011111001110111010001",
      "011101101000001001011000100101",
      "111100011111001011011111100111",
      "111110001110001101101001011100",
      "100100001110011100110111010011",
      "100111011111100111101010110001",
      "101101111011100000010110001101",
      "101000100000001101101110000001",
      "110110000110001001101000011011",
      "011000010010000011001100110000",
      "110111101001001001000100100110",
      "010011111100011001110101111010",
      "011010011111110011000011000110",
      "001101100110100110000001000010",
      "010000111101010010101000011010",
      "101111010001000101001100011000",
      "111110100101000110001001001101",
      "101101011010011110111110011111",
      "000110001010011101111101001000",
      "001110111110111001010011101011",
      "100100110010111011011100101000",
      "110110010001000100100000101110",
      "100001111101101110111011011101",
      "010101101111101001110000110110",
      "110011110111101000100100000000",
      "001111010100011001010000000001",
      "101010101110101011000011010001",
      "000110100011011110010110111101",
      "110110010001011001001011101000",
      "011001010011111001111001011101",
      "110101110011110111000000011100",
      "101001011100011111110110001010",
      "111000100100011000010100011110",
      "010100011110001101000101100011",
      "110001010000001001000101111100",
      "001000010010000010110100111111",
      "111000100011010011111100000101",
      "111111101011000110010011111011",
      "000101010001010101001101010000",
      "101011110011100101010111001110",
      "100011111101011111011101001001",
      "010110000101001110011011000000",
      "100010000100010010010111011000",
      "000100000001100111110010010110",
      "101110010110000111100001011001",
      "011001100011111001100000001001",
      "001001110101000100111110101000",
      "110100011100000011101010010111",
      "010010110001101110001100001010",
      "011100110001101011110101010011",
      "010111001000100011110110010011",
      "011000000001110111011010110001",
      "001101000101100000010110100110",
      "110001001110110100100111101010",
      "110011011001110000001000011111",
      "101111001100011100010001101111",
      "000101111101100110111011100000",
      "101010010000101111101001000001",
      "110010110110100110110100100001",
      "110101000001110000110101111111",
      "100001011010000100001100110111",
      "110010101100100111000001010110",
      "000011001101100111010101110101",
      "000001100000001001010110011010",
      "111100111010000000011000101000",
      "010110101100011011010000100101",
      "111011001100100010001001000010",
      "000110110000110011001101111001",
      "001111110111011101100000010010",
      "100001011101101100001000110111",
      "100100001100011011111101001100",
      "001101110111110001100110011110",
      "111100011111101101010100011001",
      "101101110111101010000101001001",
      "000011100000011110101101100011",
      "110111110011100110001101100101",
      "001000101000010001110100111110",
      "111001000001010000100111111011",
      "011011101010000000001011010010",
      "000001101100101111011000111110",
      "111001111000010000110010011000",
      "001011010011010001010000001101",
      "101001101100100111111101111110",
      "001001010111110110111000011010",
      "011100111011111000000001110010",
      "101001001000010100100001001000",
      "000000111010010000011101101001",
      "100010000110010111000101001001",
      "101100100000110101011011011010",
      "111100110100101011000010111100",
      "000111100011100010111111001001",
      "110001000001010000111101001111",
      "100101001001010000010101100110",
      "111111010001000010110111000110",
      "001110110010111000010101001111",
      "101010001011100111101111010000",
      "010101101111001101000110010101",
      "100001010111100110100000100000",
      "001100111111001011010010111011",
      "110101100111111011010000001100",
      "111011011001001110011011001110",
      "100100100000100100111111100101",
      "110110100100011101000110001111",
      "100100110110110100101110010010",
      "001010001100001000101001101011",
      "010010001001110100011001101001",
      "011101000101000101010110010100",
      "100111010111101111011001101100",
      "101100001000000001101010111111",
      "011001110110000101011100000110",
      "110110000011101101111011101110",
      "010010101111101010110110000010",
      "011000110000010001000010100001",
      "001110000110001101011111011110"
    ),
    (
      "001000100011000010110110100110",
      "000010100010000000110111100101",
      "010111111111100101001100100010",
      "001000101110101010100001011000",
      "111111011101000001001101000011",
      "001111000001101000110110100011",
      "010000110010100110000101011100",
      "101101111111101111110011010110",
      "010011000011100011000101001101",
      "010111111110100111001101000111",
      "100110100101110100011111011001",
      "001000011110011001000011000011",
      "001101000010110011011011101011",
      "101010010011100101000001010011",
      "101100111011101000100111101000",
      "110111010011111110001000110010",
      "100001000110010111110100100001",
      "010111001000011010110000110110",
      "101111001000011001111111101111",
      "100001110001010111101101101001",
      "100000100111010110111000011011",
      "001011111011011010010100010110",
      "000010101101001000100101001011",
      "001101011000011111100000001101",
      "001011010011111100101011110011",
      "010101101001101100110101111111",
      "001010100100001010100101101000",
      "011100000000110100000100001111",
      "011110110110111001101110011000",
      "101110110011100000001101001010",
      "010100110101100000001000000010",
      "010001000010011011000101111001",
      "010000100001010111010111110100",
      "101110100001010101000010111111",
      "111100110010011101111001000110",
      "101101100110011100110100001010",
      "011110110100011100100001000111",
      "111010000111101100111001111101",
      "001011001010111100100100101111",
      "110001111100010100001101011101",
      "100100100101101111010000010100",
      "001011111000010010100010110000",
      "101000000110001000101110010101",
      "011111000000000100110001101010",
      "100111001101111010100100001110",
      "000100000011010101101010011001",
      "111100000011010110101111101001",
      "100101111100010110010001101001",
      "010000000010001101111001111011",
      "010101001011001100110101110011",
      "000011010011011110100110110010",
      "000000101010100010000100011011",
      "100010101010001011110010001100",
      "000101000011010110011101110010",
      "000101001100100011011010001111",
      "010100111000110000011101111000",
      "100010101100010011000010000100",
      "111001010110010100100011100101",
      "000111110011010111001110011110",
      "000001000111010001001011000100",
      "110000101011010001000111001110",
      "111011010110001100101010100111",
      "101111001110010010011110000010",
      "001111101011001101101100010000",
      "001001110010000110010110001000",
      "111110111101101101011011100100",
      "000010101111111101101011101011",
      "111000101100101110101111111111",
      "001101000001110110110111101100",
      "011000010101001000001111100010",
      "001100010001001010011100110010",
      "010010111010011000111011101110",
      "101101111111101100100000001111",
      "000110111100011011011100110100",
      "001010110111111101110001111100",
      "011001100100110100000100110110",
      "111111011011010100011111111011",
      "110110000000100011111101010100",
      "111111000101011111100110100110",
      "101100111111100010010101001111",
      "001110000001000011011001011110",
      "011001110000011010000010100000",
      "000010010100001110100111111110",
      "100000101110010011010101010100",
      "110111001011010111011010111100",
      "010111000111000110101110111111",
      "110000011101011110000110011011",
      "110101101110001010010110111101",
      "000101011000011010110101010010",
      "100100100000100010100000011100",
      "101011001001100111010011000110",
      "110111110011011000001011011001",
      "111000001010111111101010110010",
      "111000111010011011001110100111",
      "100011110111011110110100100010",
      "010101001001000010101110011010",
      "101100111100101101011110100001",
      "101011110111111010000111100100",
      "011010010101010110110001101100",
      "011000010000100010001100100111",
      "111100001111001101100111111110",
      "110011010101100100111000100010",
      "111100101100110101010000001001",
      "101111101011001101010011111111",
      "100010111101000000110101101000",
      "101111000010110111100010010011",
      "010111000000110100110101010000",
      "011011110000011100001101110000",
      "000011011111111100110110000011",
      "011110100101100111001111101011",
      "110111111100000001110000001100",
      "011100010110011011101110101110",
      "100000000011111000001111101001",
      "100111100011111101111011010000",
      "011010000001010111101110001001",
      "101011110110110100011011100101",
      "100000100110100111001011010101",
      "111000010011000001111011010011",
      "011010001000010000011111110111",
      "010100001110100011110101000100",
      "010101100000111001011100111011",
      "000000100100011011001110001111",
      "111100011101001001010110101101",
      "001111110101011101101001001010",
      "000100111001111010010010011010",
      "001001000011001100111100100000",
      "110110110000010001001110010101",
      "010011101111110010100010001000",
      "101100000011100110111111101101",
      "110111001000010111011011000110",
      "100100011001000111011100011001",
      "110000111101000000111011100111",
      "101100010000101001101000101010",
      "001011111011110100001010101110",
      "011000010110010001101110111010",
      "100011100100001000101011011111",
      "001011110101001110011100001110",
      "011011100010100100010110001000",
      "110000001101010101011101011111",
      "100110010010110111001100010001",
      "010011111101111110011101110000",
      "111010010000110100110001110100",
      "000011100101100111110001100100",
      "000101011010101100011111010110",
      "010011011000100010011010110100",
      "100110110001011001110110111111",
      "011010100110011110000011100110",
      "111011111000010110011011000011",
      "110100111000110010011010000111",
      "100010011110110111100010010101",
      "010100010101111000010001001100",
      "010110010111110001001100001000",
      "011101101010011011100111001010",
      "010101111101000011101011010000",
      "111011101110100011000110111100",
      "101010100100010000110100100000",
      "011001010000101110010000101110",
      "001111010001100001010001011111",
      "010110010111001001110001100011",
      "100110111001101001111000000001",
      "011011010111111100011010010010",
      "111001001010011010111110000011",
      "110100000010000111101110011000",
      "010010010111100101001100011011",
      "100011010101111010000000100011",
      "011111110001100100010001110010",
      "100000010010111001101010001011",
      "101011100001100101001011111010",
      "100001000100001100000101000010",
      "010100010001000111000100101110",
      "011010000010000100000111111001",
      "011010110110100101111100100011",
      "011100111111010101001101000111",
      "000011101011001101111111000001",
      "000010101101001010011010111111",
      "111111011001100100100111110111",
      "001010111110100101001000111011",
      "010001101110110100111010011011",
      "010100100010000111011101110010",
      "011000000100110001011010111000",
      "110111011001111101111011101101",
      "101100011100011101011110001111",
      "000101000100110001100011001000",
      "000010011101000100000110000111",
      "000101010110111010110000101011",
      "101010010101001101100011110101",
      "111100001011100110000000001111",
      "110110111101001011000001101110",
      "101100101001101101010001101110",
      "011110010010010000100000001000",
      "101110001000000010110110001001",
      "000111011100010010011111101011",
      "010010111111010001011100001011",
      "000001001111110101101010110111",
      "101101000000110011010001011111",
      "000011101110101101111010101101",
      "111100001001000010010111101100",
      "010010101110000000101110111001",
      "111011011010101101101100000111",
      "001010101000001001111100111010",
      "101001000110010000010000100101",
      "011000110000101001110101111100",
      "101000111100110001110001110101",
      "000001000101001001110101001001",
      "110111111000001001111101101000",
      "111000011100001001101011100011",
      "000100001101111101101000101000",
      "010010111111101110110100100111",
      "110011011001010011101011100110",
      "101100010111111111101011011110",
      "011011000010000001110100010111",
      "010110010011101010101111100011",
      "011110100000010111011111110100",
      "111100100111001011001101110101",
      "111110010011011100110101101011",
      "000001100010010010011010111011",
      "001010001000011101100110000111",
      "010010000100100100001111011100",
      "010101000001011011010100000001",
      "111100111010111000000111010001",
      "000111110000100001111111100000",
      "100110110110011001110100010010",
      "111110010011011110111101010110",
      "011111001110101111000101101101",
      "101011000100011100010111001100",
      "100111000010011000010101001100"
    ),
    (
      "000011100000111001100000100000",
      "111100000001101110110000011100",
      "011101001000010101010010101101",
      "001010111101000101101001010011",
      "010101110111011111111000111001",
      "011101000011000100011010000010",
      "000001110010101000111100000100",
      "101101110101110011111100010001",
      "011101111001100011000000001110",
      "101110101011001010001110010111",
      "110100110110001001101001101101",
      "101001010010110100100100110001",
      "001111111111111111110111011100",
      "111010111100001100001111001101",
      "000000100010100001010111110101",
      "111010110111011100000001101000",
      "010011001100011010100000110010",
      "110111000011001010010000111011",
      "011001000010101001111001100000",
      "001010001000101100001100000000",
      "101001011000110000011011110110",
      "001010110010011010100010011011",
      "001000010101011001111011111010",
      "111110110000010011000011110101",
      "100000111101100011111111110101",
      "100010100101011101101100011101",
      "110010001101010101110110011010",
      "001111010100001101000111110001",
      "000111101010000101101101001100",
      "001010100110100111111100011011",
      "000100011100101010110101010010",
      "010010011101110011010010111100",
      "000110001001001101001001011010",
      "101110110111010000011001011010",
      "111101111111100111101010001100",
      "101010000100011000110110110100",
      "111010100100110000000001101110",
      "001110000100100001000000001011",
      "101111011000110101100110000011",
      "111000101010010110100001110011",
      "111101001101110110000001001011",
      "110101101110101011110010010011",
      "110110101101010011100010000101",
      "011100111100101000110110001111",
      "001110000101100101011110101000",
      "101111011101001001111000111111",
      "011101010101111110011000111101",
      "010111010100010110011011100011",
      "111011111100011110001000111101",
      "110011101100011110101100101100",
      "100000001010101111101101010010",
      "011101111010001110111001010111",
      "011010100111000100011100000010",
      "010010110001110001000001000100",
      "011100100000001000110011010110",
      "000100110111000100101010001101",
      "010101001101011101000100110010",
      "001010101100000100000010000100",
      "010100111110011010110010101010",
      "100000101000110010001010000010",
      "100101111100001100000010101000",
      "101101001000110101110110011001",
      "001101010011111100111001111000",
      "000110000111011101110100111100",
      "001011101100011001100101100010",
      "111010011011111011011110111001",
      "110000011111111101010000001110",
      "111101001001111110110100110110",
      "111011001011001011110100000000",
      "111001011001000100100000011010",
      "011100100110011011111111010100",
      "000001011000001110000000101010",
      "011110111110111101010010110011",
      "111110100111111001001001000001",
      "100000000010100100011101011110",
      "111100000000110110010011110001",
      "110110000101011111100000100011",
      "010110111011001101000100101100",
      "111001101101100101101110001010",
      "001110101010011001101110110010",
      "101001110110101010111010100100",
      "111011100100101100101110110110",
      "101111001101010001001010000101",
      "100001011000001000101001101111",
      "011100000110101101010001100010",
      "010110001001010110101110101101",
      "111100011101101010100010111001",
      "011110111100011000101110110010",
      "001110010010110101001011010101",
      "001101000101111001001101010001",
      "000010001110001111000100000000",
      "011100101111010010110101011010",
      "100000001011110100011110101001",
      "111001110101011101101001011000",
      "100101010111111111010000110011",
      "110010101101001111100000100100",
      "111110100010100101110010100111",
      "011011000111100000001000001100",
      "100001001011010101110011100110",
      "101110000110101001110010001111",
      "000000111000011011111111111000",
      "001110000001110011010000110100",
      "101100101011110101101111101011",
      "100001001000001101000111000011",
      "001010011011010010101110111001",
      "111010110100110101101001001010",
      "010010011000111100010010100101",
      "100010001001001001100110111100",
      "110011001100101011001011010111",
      "101100110001111001000001110000",
      "000100110111000110111100100100",
      "110011000001110001100100000010",
      "111101110001011110101111101010",
      "001011111110001001111010111100",
      "111010100000100000110110111110",
      "000000010101110100111001000101",
      "100011000111100111011101111001",
      "110001111111101110000010101101",
      "010000000010100000111011101011",
      "000100101101110000011100000011",
      "011101111001001011101110011100",
      "011000011101010110010110001110",
      "000111111000011001011011001101",
      "100001001010010011011100010110",
      "011001011011101110111001001110",
      "011011100110011111000011010100",
      "110100011110011010101101100111",
      "110110100000001111110011110110",
      "001001011100011111101101001100",
      "011110011111110011000101000110",
      "001101101011111101010111000101",
      "111101010111000111101101110010",
      "001001011011011011110001110100",
      "001000101111011001011110001100",
      "100101011101000001001111111011",
      "100111000000010100111101011001",
      "011000111010100100010000100101",
      "100111010111111110011101111110",
      "111011000111010011100111111001",
      "011101000011010101101011111010",
      "100000100100111100001010011000",
      "011011111010100001110000011101",
      "100100000101101101111001111000",
      "001001010000111000010000100100",
      "001100001001101000100101001001",
      "110000010000101111001011011110",
      "110100000100111010000000100010",
      "111000001000110110001000010110",
      "010001010111110011101100110111",
      "100011101110010111011101111010",
      "100111110001101111101111001001",
      "110110100010111111110101101110",
      "010111100001001000100001111011",
      "010110111101010111010101111010",
      "010000010011000100010111011000",
      "100101000110001000001011011011",
      "010000001100111010001110101111",
      "001011100010011001101100010001",
      "110110101001000101011100100010",
      "110001010011010101010001000010",
      "010001010101100000001100101101",
      "011010100001111111111101001100",
      "100011000000001000101110011110",
      "000111101000110101100100011000",
      "000011011011000111000100010101",
      "100101001010010100110000011100",
      "111000111101010100010001010110",
      "100011010111111001111111011100",
      "010101000111010010110111101001",
      "111101100110100111011001011001",
      "000001110010110000101100011000",
      "100011010110101011111011111011",
      "110110110100111101011110000010",
      "010110100111110110000001001011",
      "100010110100110101001101011000",
      "010100000011000110110101011110",
      "001110100110111001110010110010",
      "010111100100110010010110001110",
      "100000111001111010011010100100",
      "000001100110010100011000100100",
      "111011101110111110001110011111",
      "011011101101111100111011000010",
      "011000101100111000110011110010",
      "100011100100101100101000000000",
      "000101100000100100011001111011",
      "010101100110000101111100111111",
      "000001111001000110001000000001",
      "100110110100100011110111111010",
      "100001111011000100111000001001",
      "100101011011011111011011010000",
      "001110111000101101111100001110",
      "100101100001100100101000111111",
      "111110001110100101011000101111",
      "000110110001000010010000100110",
      "011011110000001101110110100001",
      "001100110010110100011101111001",
      "010100000110111100011101001001",
      "001101111010001010110001001001",
      "111101110000010011011000111101",
      "111011111111000100011110011110",
      "000101111110001011000110110011",
      "111100000011011010010000101000",
      "011010110111010001000010111110",
      "110001100101011111111000010010",
      "111010101001101111010010101010",
      "010001101000010010110010100111",
      "000010011011000100111111011101",
      "000010100001011000000001001001",
      "000011000010000011111100001001",
      "001101100101011011110010001111",
      "011011011101110101011101111101",
      "011000111111010101100010100100",
      "011011000111010111000100100110",
      "111100011011101000110000001011",
      "101011011000101111110111000111",
      "101011111010000100110010110000",
      "110101110010101101010101110111",
      "010001110000110001111101001101",
      "001110110011110011101101110101",
      "010001001011111010111001001111",
      "101001010000000001001001101100",
      "111111011001011011100101111100",
      "110100110000011110001010110101",
      "100100110001001000100000100110",
      "000111111100000101000001111011",
      "110101010001001011101000100010"
    ),
    (
      "110110110010011000101101110010",
      "101111111110110011011010101101",
      "011110101000101000101000011010",
      "001101100000000010110111011100",
      "101111011011010000011000001000",
      "101110011011101010001110110111",
      "111011101010010010010110010001",
      "001000101000011111010110110000",
      "000100110011010110110000000010",
      "011000111000011110001010010011",
      "000111000110010111010101000111",
      "000100100101010001001100010001",
      "000000010111101100101111011000",
      "111011000111010011010011111010",
      "111110010110011000111111100110",
      "000011100011111000110001110100",
      "010011011000000001100100011010",
      "001100010101001111001000001110",
      "011000011011110100101100111100",
      "000101101110001011011101100001",
      "011111000100010111011100001001",
      "110000000010101011101010001100",
      "000100000010001011100110110111",
      "011010011010101011111001111011",
      "010010011100100100101101111101",
      "110000101000001100111100000110",
      "010111001000101010001100110000",
      "100100111000000110011010001100",
      "100010110000100100010001001111",
      "101111110010011010100111101111",
      "011100100011101000011100101010",
      "000110100011111000010000010111",
      "101001101000101001101001010100",
      "011101001101000101101000101111",
      "110000010010100110011111010100",
      "110111100010000000001110111011",
      "101010010101101001011010111011",
      "110001000011000111010110000000",
      "001001111101010101000010101100",
      "100011110001001100011001100111",
      "110001100001111111111001110010",
      "011001101000101101000001010101",
      "110000011001100110111011111100",
      "010101001001001100011010100111",
      "101010101111001110001110111110",
      "111001110100100101011001010100",
      "001101011001000100010101101010",
      "111001010101000011110101000000",
      "001110100110000100001111110100",
      "000100111010110010101100011100",
      "111101001110000101100010001001",
      "000000001011100110101100000111",
      "011001001001111010001101111111",
      "100101100111100100100111110110",
      "010101011000111000010111011011",
      "011010100000101101010000111000",
      "010101100110100101000100001100",
      "010010010001101110001011001111",
      "010000100011100101110010010110",
      "000001110010100011100100000100",
      "000100101100001110111011010110",
      "010110111001000001010001111010",
      "101111101111001010100110001101",
      "000001000100101100000010010001",
      "011111110001101000001111101011",
      "001010110110110011110011010100",
      "101100111010100110111011011001",
      "001011101001110111010110101010",
      "000000010010011011101000000111",
      "100100101111000000001001111101",
      "100111101110000001111111001101",
      "000111010011100100001011101111",
      "101111101010111000111000111000",
      "001111001011110011000100101001",
      "010101111100011101110011001000",
      "011000000100100110111111011010",
      "000001000101001010001110001110",
      "000111110101000110000010101010",
      "111111000011101100110010111111",
      "001100100111100011001101000000",
      "110001011001010100000111100110",
      "011110000000011100110000110011",
      "110001001000000010010100111011",
      "110000100111111001101100010010",
      "010001010101111110010010011111",
      "101111001100110101010111010010",
      "001100000100110001001110101011",
      "000001101100001001000110100011",
      "000101011000001101100110000011",
      "010101000111111000110010111111",
      "010010000000000010100000111110",
      "110110110101000000110011011110",
      "110001111110010100011100011001",
      "100010111111001101111111100110",
      "010011100111001110111110000001",
      "100001110100011110010010110000",
      "100010011010000001101110111111",
      "101011001011011001010011010111",
      "111010011110010110010111101010",
      "111000011011111101011011011010",
      "011000001000011000101110000010",
      "110010010011101011010111010111",
      "000110010110011001111010010001",
      "100000010100011011101101110010",
      "110110110100001100001110101000",
      "111001100110111101000110011000",
      "101011001100000110111100011011",
      "010010101011001110100110000010",
      "010011100011100111101110100000",
      "010011010111110100001100001010",
      "101111101000011100001111011111",
      "100000111100101010101101101011",
      "000000101111111000001010100001",
      "111111000011000010110101110101",
      "111010000000100100101101001011",
      "110000010111000101101111011011",
      "101000010011101101111011110100",
      "001010001111111110000111101100",
      "010010011101101001001101100001",
      "111101100100100101101111110011",
      "011011010001101101111000101000",
      "000011111001000010001101001000",
      "001000010000101100101011111011",
      "001110011001000000000110100011",
      "111001101001011110110001110010",
      "011011110110010000110101000100",
      "100110001000011111110101000111",
      "110011000100110011000110001111",
      "001000111111101000111000001101",
      "000000011100101010100111110001",
      "110010000011100110010111101111",
      "101100111110001111110010111010",
      "010101101101110010101111001000",
      "100111000110000011110111001000",
      "110110001100111111100000111001",
      "011000001011111101010111010101",
      "100010111100011000000000010100",
      "101001010001110101101111010111",
      "101011110100000010100110001110",
      "100110000111001111110010101101",
      "000011100111001101101010000001",
      "011010001100111101111101111110",
      "111000101111001101010010100101",
      "110000000111101001101001000000",
      "010000101110010011100000111111",
      "100000100100111100111010010010",
      "101011101101110110100010011100",
      "110110111011100101000110011111",
      "000011101000110100000110000001",
      "100111010000001111011011000100",
      "011111000101100000000111110011",
      "000001110001110101110000011011",
      "011111000011111101011100011000",
      "100010010100110111101101111101",
      "001110000011111001111001001110",
      "110001011100010110000000100110",
      "111000011010011101001111101000",
      "000110101010000110001101110110",
      "101101111101001101100111100111",
      "110101100110111010011000111111",
      "000001101010101001011010011101",
      "110011011101111111011111100001",
      "110111101111010100011001101100",
      "001110001001010100100111111101",
      "101000100010111110100111011111",
      "100011110111010101001010100111",
      "101111101100111001100101111110",
      "011010011110101000110101100101",
      "010111100001000100011011100101",
      "010111101111110000011111110011",
      "110011100010110000100000010010",
      "001100111100100101110100011000",
      "001001011000111101100000100011",
      "100001010010111110011100100000",
      "101000000010010011010010001011",
      "100101101000001111000010110111",
      "000001111111011011001000011010",
      "100011010111110111110100110110",
      "100000010110011011001110010111",
      "110010100101111010000111000110",
      "000000010111000010100000000011",
      "101011001010001110101010011010",
      "110110101100100001001100100010",
      "000100000111100010111010001111",
      "101100010110101111111110110101",
      "011101011111001010001000010101",
      "001110011001001000001010110000",
      "101101101110000101001100100001",
      "101010010110101101010111101010",
      "111000111001110010111110011110",
      "011011011011110001001100101001",
      "110111001101001101111101011000",
      "101110100100101111010010101001",
      "101011101011100100110110001011",
      "000000000000010000000010111011",
      "110110110110101010000110010001",
      "101111001011001101000011100110",
      "111011101101100101001011000110",
      "001000101001010001100001011110",
      "101100010111001100100010100111",
      "010010110001010011111111000011",
      "111101001010001111001010011010",
      "110001000101011110011111101111",
      "111011011101111000001001001000",
      "101011101010100100110010110101",
      "010010011101001110110000001011",
      "111110000011000101000011011000",
      "110111011110010011011101110111",
      "110101100100001011010100110000",
      "100001010001001110110111110001",
      "101101010010101111100000111101",
      "011001100001011001010101110010",
      "010011011100111011111000101000",
      "010111011101000011011011010001",
      "010100101000011110111010101011",
      "001111101111100001000011010001",
      "110111111101111110011110001011",
      "100011001101111111100110101100",
      "101110001100100000011001110000",
      "011010001111111001011111000011",
      "111111001000111000010110011001",
      "110111111010000110100101111010",
      "110010010111011011011100100111",
      "101101101111001011010110011001",
      "000010110011101101101111011000",
      "011011111110000000100110000000"
    ),
    (
      "110010010111101000111100100101",
      "001010110110011000010110001110",
      "010001111110011110101101011111",
      "011111001011011010111111000000",
      "001111000001110111111111010000",
      "111010110110100101111001111010",
      "001011001001111010011010110000",
      "011111001100111100000000010010",
      "000110001101001101000010100001",
      "001100111000110011111101111101",
      "101100110011101100001010101101",
      "011010101110010100010010110011",
      "100010111001110000100001100011",
      "101010011101111011001001101101",
      "111110100010011000011000011000",
      "001111101010000110111000010101",
      "111100011000000010101111101001",
      "101101100110000010111100000111",
      "011000010011001101100011111011",
      "110011000110000000111010000001",
      "100110110001100101010001011010",
      "000000110111111100000010110000",
      "010011001110110100010110100000",
      "111100011001100111011110011010",
      "000100110111010000101010011011",
      "100111100100010100001000101111",
      "000000010011011100101101110101",
      "101000111100101111011101000101",
      "001110010110110010111100011100",
      "001101101001101110000111011001",
      "111011100000100011001110111000",
      "100011100000110100111110101110",
      "001110110100011110000101000001",
      "001111011010101001000000001111",
      "010011101101100101001011001110",
      "100100000011100101010011011010",
      "101110000111111000101001000010",
      "001111011010001010101110001110",
      "111110001001101011110110011101",
      "111100111011100101011100100010",
      "101010110100010000100010010000",
      "010011011001000110111100100010",
      "100000110000010011011000110110",
      "010111101100111000001001011111",
      "110001000011000100010011000110",
      "001110011111001111001000110010",
      "011100110000110111000110111100",
      "100111011000101101001110000011",
      "100100100111111111010001111100",
      "110001110010001111110000111110",
      "011011110101001100000110111010",
      "100000111100011100100010111010",
      "100110000100001111110010010100",
      "001000101011100010110100010111",
      "011001111011001101011111000111",
      "001001100000111101111000010100",
      "100001100100100001010000110101",
      "110110000011011011110001011001",
      "001010000101100110001110101011",
      "001000000110101111001000010111",
      "011000110001011011010001110011",
      "000101110110000111110011101000",
      "000000100011001000010110110010",
      "110010010110001111100101000001",
      "000000011100100100100010010011",
      "000101000111110110111010111111",
      "110101001111011000000101101100",
      "111000001100111010011000100110",
      "000111010011010111101010000100",
      "101111110010110100100101000011",
      "011111111101100010100110111100",
      "000100101110101111011110111111",
      "101011001100001101000010000010",
      "001111001010000111000111101001",
      "101101011101110001000100100101",
      "000100101011110001011011001100",
      "010001000110001100000000100011",
      "000101011010111101111100000000",
      "001100110001101000111110101110",
      "100000000111000001001001100011",
      "001100011111011011110110011000",
      "100001010101000010001000111010",
      "011101101001000000011000100001",
      "101011010110000110010000000001",
      "101110111001110010011001101001",
      "001111000111100001010101000010",
      "010000101100000000110111010001",
      "100010010110111011011001101011",
      "010101011101000000111000111000",
      "110000110111010100111111111001",
      "010001000110001000100111100000",
      "110001010111010101111010101100",
      "101111100110011001100000001000",
      "100001001000001111011110000000",
      "011101011001101010111101001100",
      "010110010010010001001101001010",
      "001011111100100010001001101000",
      "101000011000100101111010000101",
      "011111001000000101011011111011",
      "000100000000011000111000010111",
      "111000010111101010001001101111",
      "000000000111000100110111111001",
      "001110110010000110010010001011",
      "110001001111000101010010101000",
      "001100110000110110101011100100",
      "011100001111010010011010011011",
      "111111111100100011000011010101",
      "011100110111100010001001110101",
      "001111011011001110011010001111",
      "000101110000011000111111110111",
      "110110010111010010100101011000",
      "101100101100001111010010101111",
      "001100000100000110000010000000",
      "011111101011110110001011001000",
      "111110011000110110110010101000",
      "011011101100010001000000101101",
      "001001101010011000001100010000",
      "111000010011101111100010111110",
      "011001101010010010100000010111",
      "001011001000001011000110010101",
      "100010100110111011010010011011",
      "101101100100000110110100011100",
      "100110000000001011101000011000",
      "001111110000011001100001110110",
      "110110100111001110011001010001",
      "011011001111011100011000000010",
      "100000000110011111011000110100",
      "001000011000011110111101101110",
      "111100001010111101000101100101",
      "101001010111001111010110101001",
      "101110111011101010000101100010",
      "111110100100010001011110101100",
      "010100001001101110011011001101",
      "110010100110111110100011011110",
      "000100101000101011110110011110",
      "110111000101100011100010000010",
      "111011101001111101101100100111",
      "111110000001100111001111001111",
      "010001010101101101011010100110",
      "111111111010001001110101001101",
      "000000110011011001010110110111",
      "110111001000101110100010001011",
      "010001101001111001101011011010",
      "110111101111010110101010001001",
      "010100100010101101010100111000",
      "001111101110000100110100010100",
      "111001000100100011010001011100",
      "000101101010000111111101100011",
      "001111000011111001000010101101",
      "111100100010010101010111100100",
      "000011100110011100010111100001",
      "100111000001111000111100001000",
      "111100111011110111100110110110",
      "111110011111100010000000001001",
      "100111000100100011001110111000",
      "001010011000111001100010100000",
      "000011101000010001000101000001",
      "100001010011010101110001101011",
      "100011010011110000101010010101",
      "100110100011000011011100101101",
      "010101100100111110100110011101",
      "101011111000010111011101000000",
      "111010011011010100000100101110",
      "010101101000111101101111010110",
      "010011110111010101000001110111",
      "110010001011111011010011011111",
      "000010110011001110111101110011",
      "010111110000110010000110110111",
      "001110000000110110111001011110",
      "001111010110101110000010101001",
      "010111011010001100100111000001",
      "110000001011011010001010001100",
      "110111011001111001111111000000",
      "110000100111100110001110001110",
      "000001011101100011110011101110",
      "100010000100110101101010101100",
      "011100001011001011110110000100",
      "000110010001000111001001111001",
      "000011111001001111010001010110",
      "010001010101110101111000110111",
      "100010111110111100101001110010",
      "001000010100100101110110000001",
      "010111011100110011010110011100",
      "111011111010011111010000001111",
      "111011101000110000000110011000",
      "111000010110111000000111000011",
      "011101111100110001001100110100",
      "001001110010111001010010111110",
      "110101101010011010010111010010",
      "111100001000000000111000001001",
      "010011110011100111010101011110",
      "110010001011011100110001011001",
      "101110011010101000010010100000",
      "001111010111101011011100000000",
      "001111100100000001111011010100",
      "011000011110011010111000111000",
      "011010000101110010001011010111",
      "001110110111010011000011100111",
      "001001011110101011111001111101",
      "101010111110000101001000011001",
      "000010010110101010001011101010",
      "000001000110111101101011000111",
      "000011001011110111111100100110",
      "111001111111011100100001110010",
      "001001100100111111010110111000",
      "111100101000111100000011111011",
      "100000000000010100110000010101",
      "110001011000110011010101111100",
      "100110101101010011101100011010",
      "110110010100011010110000101100",
      "010001010001010001010010000010",
      "010001110001100001101110001101",
      "110101010001111000100011111111",
      "100001010001100111001011011011",
      "001001000111011011000000010010",
      "001110010110101111100000000010",
      "010001001000110000010001011010",
      "101100001101001000111010000110",
      "111111000111111001000000111000",
      "110111010101101110000000100110",
      "110000011011000010101011010100",
      "011101101010010111010111100110",
      "000100111110100111100100101000",
      "101100011111001010110010100000",
      "111011110000101100110010001000",
      "010101100111111011010110010000"
    ),
    (
      "110011011111011001100100000001",
      "010111011101000101101010011011",
      "110101011110111010000110110101",
      "111110111000111101000011000010",
      "110100111011001010011010001110",
      "010101111000011100001011110100",
      "100100010110011011100110110010",
      "011110001001111110110110011110",
      "000000111000010100011111101111",
      "001110010100111101011111100001",
      "000111011111111110110110110001",
      "101100111110101000101011010000",
      "011011011101010100001001000000",
      "111001110100000101111001100111",
      "110101100000111010110111010011",
      "011010101010111001101111100110",
      "111111110101100001011101110010",
      "010011110111001111010110111100",
      "100100001001011110101000001111",
      "100001010110010010101100011010",
      "001111101000001110100110000101",
      "111010010111100111011010000101",
      "100011110000101010101001000010",
      "001011100010100011110100100100",
      "100110011011000110100000011001",
      "001001010011101011100110011010",
      "101000010110001011010010010010",
      "000101000000010111000101110100",
      "010111111000011111110101110101",
      "111001100011011011001010110111",
      "011000111110000100000101000001",
      "111001011011111110111100010110",
      "110011111111110110010110011101",
      "101011001101000000100000110100",
      "010000010001101110000110110101",
      "000101011101100110110010111000",
      "100011001000100010111111001101",
      "111011111011100101001110110111",
      "011101000101101111101001100011",
      "110010100000110110101110001100",
      "110100001110010000010000010001",
      "110011110000001111001011101011",
      "101001011111011010010100011100",
      "000011001110100000111000111101",
      "101011001010110011101111011110",
      "000011000100010001101110110111",
      "110110111100110101101000110010",
      "011011111101101001000000100000",
      "111001000111001011011011101001",
      "101110101100100110000011111100",
      "001100001011011100101010001100",
      "111101111100000001100101110011",
      "100100100101111100111111111010",
      "101101000101111100110111001111",
      "000011111101010010111000001000",
      "111110100110110001111110001001",
      "010011100110101101111010001111",
      "101101101111110110011101111011",
      "011100011011010111100100001101",
      "101000110000111010010100010001",
      "000000100010110010110010111110",
      "000010001010110011100101000100",
      "100011011000000111001001111001",
      "101011000110101111001000100100",
      "000000000101100010011101010001",
      "011010101011011110110110101010",
      "110001101000101000100111101110",
      "110101110111001011110001001101",
      "110011001111101101001011101101",
      "001110001001100100011001000011",
      "000101011010100100000010111101",
      "000110001100010100010001111000",
      "001100111110110001000011010011",
      "100011100001011010010110110100",
      "100111010111110111110000110100",
      "001001110111101010110011101010",
      "011010001101100010111000001101",
      "100101101110001010101101110000",
      "100011111111110111100000111001",
      "100000100000110001001100110011",
      "001101111100111000000111000101",
      "111010001111111011110001000111",
      "111100101011011110001011100101",
      "000101001000100110100001010111",
      "110001011000111001100001000011",
      "101000110101011101110110010110",
      "011111110100001010101110101010",
      "111000010001010001001110001011",
      "011110010101100010110101100101",
      "011001010011111010101001111111",
      "101111000101101000100110111100",
      "000000100111101010011110001001",
      "100101111000011010101010010011",
      "111100110100110010100100101111",
      "011011000110011001101111100001",
      "110001100000011100111111010111",
      "011111000100110001010111001110",
      "100000100011011110101001010011",
      "000000011000010010100111110000",
      "001101110011100111110011000100",
      "010101001000110001100111101000",
      "001100101010111010000011000101",
      "110111011110010101000011101000",
      "111000110110101011111100001101",
      "000101001010011101100100111111",
      "111001010111100110011110110101",
      "101111100110100100110011001101",
      "111001100001101011111011100010",
      "010111000011001001101100101101",
      "111010001011000000000001001011",
      "001011101000000110110010101010",
      "110010111011111111011110111001",
      "111101110111101010011100101011",
      "110101010001101110011011011001",
      "110010111100101110001100000100",
      "101101111111011000011011001111",
      "011111011100001011010000001110",
      "000110101001011010001010011100",
      "110011101100010110101001100010",
      "010011011010001110010001101101",
      "011010010101110111101000110101",
      "010000100010010010110010000110",
      "111000000111001001101010100111",
      "010000110110100111010010000000",
      "011010110110100010010001010000",
      "000111011011111001110111010000",
      "011000010001011110100010000101",
      "000100011010011010011001100010",
      "011100100011100001111011000000",
      "101110111000011101100000111101",
      "011110001101101010001010001111",
      "101100111110001011000001011000",
      "000011001011011111101100111001",
      "000000100101000101011100101011",
      "000111101100111100101111010000",
      "000001100000111000101000001001",
      "111100001010101100011101010001",
      "101101111001110100000011010000",
      "101111001000110001000111010011",
      "011001100000011101010111000110",
      "011111101000001011001110000010",
      "000101110111100110111100001011",
      "011111111010000110001011100101",
      "001101011110100000001000001000",
      "110100110011000101011001100110",
      "000000010111011111010111001001",
      "101011101010101011000011111110",
      "101010110100110101101100011010",
      "110110101000110001101010101001",
      "010100011001110001000110011110",
      "100110010011110111101101010111",
      "010000001011100010000101110010",
      "010101001001011010011110100100",
      "110100010111100001011100011110",
      "101010010001111010010000011111",
      "110111100110000000000001110111",
      "001011011101110000100001001010",
      "100010001011111111010110110110",
      "010101000100010100101010111110",
      "011010001101110011000001010001",
      "010000101101000000110101111010",
      "011000110111000001000111011010",
      "100110100111100100001000111010",
      "111011101100010100100110001110",
      "011010111010001101011011110001",
      "001110000111001111101110111001",
      "010010100001101001101011001000",
      "001000110011010011001100010111",
      "101110110110111110101001000011",
      "011111100111000101001100010111",
      "101101011011100000010110100011",
      "101001010111000010010111010011",
      "101001010011101111111110000101",
      "011110000101000010111101011001",
      "001001000010110000110010101011",
      "001110111000001111001010100111",
      "000010110100010011100100111101",
      "100100011011100011011101100110",
      "100010100001100101001001101101",
      "001100100001110110011110110111",
      "110010011101100111000011011110",
      "110011111100110100100100011011",
      "011100010011111100111110000101",
      "111011111100001011000001100011",
      "111011110000101001001010011000",
      "001011111100101011011011100111",
      "101011001000101101010100010100",
      "100010011111101000111001001100",
      "000100001110100111110110001001",
      "111101001101110011010010011000",
      "110101100000000011000000110100",
      "011110111110101000110100011111",
      "001011101000100011011101101111",
      "110011000000101111010100101001",
      "101011010010001111001010101010",
      "101011100111010011111001011100",
      "100011101011101011101000111101",
      "001001001111000101111000100111",
      "110011110010100100000011100000",
      "000110111000000110110011111110",
      "101011110001100101001010011000",
      "001110000101001000001000111000",
      "101100100011000110110101101110",
      "110111110111001011111011001101",
      "011011010010000000110111110000",
      "010010010010000010010100110101",
      "011000111110101101111111110010",
      "000100110111000001010010000010",
      "011010010110011111100111010101",
      "011100000111011000110100010110",
      "101001001111000101001010001111",
      "110111001110111110000011010000",
      "111101100110000011010011111111",
      "010010011011100111101000100010",
      "110101011000000000011000001110",
      "011111110100010100100100111001",
      "101101110000011001110001001011",
      "110010111100100101101100011000",
      "101011000000000101111010100011",
      "111111010010101110110001010000",
      "011101000111111001010111101100",
      "101011000101101110010101111000",
      "011111100101010000010000100101",
      "011011011110110100111111001011",
      "010011101010010110000011011110",
      "111111101001110011000111111110"
    ),
    (
      "111000110100100010001111111110",
      "100000000001111110011000110111",
      "100000110001000000111001111101",
      "011010111111010111110010001011",
      "001110100101001011101010101111",
      "011011000100110011010111101100",
      "100011101001010100001000011110",
      "100011100010100001011011111010",
      "101110011101100010001011010000",
      "100001011101110010111011110101",
      "110001001101101111101000011110",
      "011011000101000010010011000000",
      "011001111001001000010110010100",
      "110110110110110000100011011010",
      "111100011011100110101011000001",
      "100011110010101010011111010110",
      "010010100000000111000000011000",
      "101000110010001100110101100111",
      "111100110000001000111000011110",
      "001110000010111011110010001001",
      "101001111111111010010110011110",
      "001000001011101110010111010101",
      "000010100000010110111000000110",
      "010000011010011011100010000110",
      "110000100111011111101101011001",
      "110110110010100010110011111000",
      "000001011011111001011000001111",
      "011100100001010100101111111011",
      "000100100001111100000000000001",
      "010110001000110110111001010111",
      "110100100011011010010111010000",
      "011001010100100011110110011111",
      "001101000110011011100101000011",
      "111011111001110000110110110111",
      "010001100010100100111110101010",
      "011001001110011001111001000001",
      "011010000000100001101011110101",
      "000110010010101000000111111100",
      "101101010101000110010001010000",
      "111100100100000111101100000010",
      "101010010011101111001010101001",
      "111001000001010100000001110011",
      "011100000110000011000101110101",
      "100010110010000110100011100011",
      "101111110111000011000101111100",
      "011000001101001101000011011000",
      "000000101101001000110110101111",
      "100111000100101001111010011011",
      "101010111000000000011101101011",
      "110111100110110010000100011110",
      "101010011100000111100001001011",
      "001010110001001010110010001101",
      "011101001011101110011001101101",
      "101110100101111111101111110001",
      "110011000100110000100110100011",
      "010011010100000010111110000101",
      "010111101111101011100111111001",
      "100111001000111111001010100101",
      "010000111011010010010011011001",
      "110110100000111100011000010110",
      "101100000111101111011110011100",
      "110110001000111010101011110100",
      "111010111101101000101101000101",
      "110000110011001111100011001100",
      "010100010000001100000001110100",
      "100101011111100001001010011111",
      "110000101011100100100111001000",
      "110010101001000111111111101010",
      "001101111000010101100010011010",
      "100011010011011001101001011111",
      "100000011110100110011000010111",
      "100000000101000010011110100100",
      "110001010010101000011010111011",
      "001000100100100101001001111100",
      "000001011110001000100011001011",
      "101111001011010101110000011110",
      "110110101100100010001001011111",
      "101101011011100111011000110110",
      "000001111100011010000001101011",
      "111000101111000011110000011110",
      "111111000001111110001111110001",
      "001000111101001101101011110111",
      "001000111011010111001011010001",
      "010111110110100110001010010010",
      "010000001110011001000011000000",
      "001101100011101011000111101110",
      "010010100100100010000000011000",
      "111100001011100100010011010011",
      "001111010101011010000011010010",
      "000101010110011100111101101111",
      "101111100100011000011110010100",
      "000111000010101111000110111000",
      "001000100000101100011110010101",
      "111000100001110010001000000111",
      "000011001001101011000110000011",
      "011101010000001111010100101000",
      "001010001110010100010010100111",
      "000001001011000010000110101111",
      "110001010010100000011110101010",
      "000111000101110101110110010101",
      "011110110011001110011010111011",
      "000111111100110011000001100001",
      "101011101101101001011100100100",
      "101000101101010110100111101011",
      "110010110001100001011001011000",
      "010111100011100000011100100101",
      "110010100100001011010001110010",
      "101000011101010001110110010011",
      "010110100011111010110110011100",
      "000100010011110100100101000111",
      "001101001010010100001100001111",
      "001111000101101001011010110100",
      "000010000101000110001100110100",
      "110101011010010110011100000010",
      "001110011001011011011010111010",
      "011111101101011101010110000101",
      "100000101000111111011101011100",
      "010001101000111000101001100110",
      "000010111011000000001101000010",
      "010001001110110100110100111111",
      "010101001111011100110100111100",
      "101001101000111011111100000100",
      "010000011100111000101011101000",
      "110111011011010011101010011110",
      "011000001111101100111010000101",
      "001001001110101011001100011100",
      "111000101010001110110101011111",
      "111001100111111011010110111111",
      "000000111001111101001110011101",
      "111110001111110000000000000001",
      "110010111000101100101001001011",
      "101110010011010011011111110111",
      "110110101110110111011001100001",
      "011011110001010011011110111101",
      "100101001111101001101000111110",
      "101010000110000110010110001111",
      "011010111001110111100110000100",
      "010110011100100010000111110101",
      "100101010111110100001100110000",
      "111010111000000001011100000011",
      "100010111010011010100101110100",
      "011000100001101001010001100100",
      "010001000111111100101000101011",
      "100110010111110110011010101001",
      "100011000000111101111011100010",
      "010101011010101100110010001000",
      "100111101000110100100110111111",
      "111110110000101100101110000000",
      "100011101111000001011100100111",
      "110001011110001100110001101100",
      "110111010011111011010101101000",
      "001011100001111110011010010100",
      "101000000111101011011111101100",
      "101101101000011101101111000000",
      "101011011110010010011110011100",
      "101000111110101010100101010001",
      "101101101001001010110000110001",
      "011111110010000011111101100100",
      "000000100110000011110101011100",
      "010010111000100011011000110000",
      "100110100011011110100101110011",
      "100111000001011000010110001001",
      "110110001010100111111011001000",
      "010001111101010011011100101000",
      "110110000000010100110100111011",
      "100111101000101101110110110111",
      "101101010110000111011001010010",
      "000100010111000011100101000101",
      "100011100111011011000001001001",
      "110101001001111100111111010011",
      "110000010010011010101011011011",
      "001010110000000111100110110110",
      "100111101111011110101001110001",
      "011010101001000010100100001000",
      "010101100101001010111111111110",
      "110000111111100101001111010110",
      "001001001011010000100100100110",
      "100111011101110000110100011001",
      "111001101000101111110111011111",
      "100011111111010111010010100000",
      "011011110010100001011101100111",
      "101110100011101001010000110101",
      "100111001100001010010110000011",
      "110110011001000100000111000110",
      "110111000010011001110011110010",
      "111011010101110110101000110101",
      "111110001111010101101101001010",
      "100110001001110111111101001011",
      "001000000000010101011011100000",
      "011111001100001110000000111111",
      "110011101101101101001100101101",
      "110100110001100111111101100100",
      "001011100101111110110001110110",
      "010001011100110011010101101111",
      "010100111000111001110001110011",
      "100101111011001110111010001001",
      "101011110100111011000111000000",
      "011101100010011000011100110110",
      "000101010110011110110100111111",
      "100000110001100011111010101000",
      "101010011101111000011001000110",
      "110001110000110110101011010101",
      "111101011101101110100100010111",
      "001100111101001110100110011001",
      "011001110111000100101000000101",
      "110011001111001001011101011011",
      "101110111100110010010100000111",
      "110110110111000010101001111001",
      "011001011010111010000100110001",
      "011000100100001111011110100110",
      "000111110011000000111011111100",
      "000001011101110101001001101111",
      "000101101100111111011110100110",
      "101000001010010000110110011111",
      "001011010101100001101000100110",
      "010111001000010101000010101000",
      "100001010001111100100101010010",
      "010010111001110001110111111101",
      "110001000010100011000110011110",
      "011101110010001110000101100011",
      "101101110011011010001101010011",
      "111011101011011010100111010011",
      "110011100110101101000000101110",
      "101001001100001011010001000010",
      "010011100110001101010111010100",
      "100000110101000010011100010000"
    ),
    (
      "000010101011011111001110111001",
      "010111010001110000000011010011",
      "100100001000101110001101010001",
      "010000010010000101100101110011",
      "010010001001011110000111111101",
      "111011101100101101110100101011",
      "000101000101011000111110001000",
      "111001101111110000111010110010",
      "110100110101011101000110110011",
      "101001101101010110000110010100",
      "000100010010110001100000011110",
      "010000000111111110100001101100",
      "110001111000101001001000000110",
      "111100010100001101111010101001",
      "011000001101111001010010100010",
      "001001110011100100100101111101",
      "101001011110010111010011100011",
      "110101011010100001101000010001",
      "111110010111101111110001111111",
      "110110111111000010010101101111",
      "100010000001101100111101001001",
      "010110101111100011010111011100",
      "101101101100011101000111101111",
      "101011101100011110001010010010",
      "110000100010011101000101110000",
      "001011001111110101110100101011",
      "011111101111101001000011101111",
      "010101110011110101100111101110",
      "001011001111100110001010011010",
      "010101100111111101001011100100",
      "001010011000011011101100111101",
      "011010101100111011010001000011",
      "010100000010101001001011010010",
      "011101000010110100101110101110",
      "110010111010100001100101110000",
      "110110010110100110001001100100",
      "011010100011101000011110100001",
      "010100101110000001010010010001",
      "011011001001110110001101110001",
      "110111011011110100000010011001",
      "011101011011011101100101010101",
      "001000011001110111010010101110",
      "100100011000101110000011010000",
      "011000011101110101110110100111",
      "010010010010010010101011011110",
      "100010110010110100110111111101",
      "001010110111110100111111101000",
      "010101111100111110101010011010",
      "111010000110000101111010101011",
      "110111011101011011000011101011",
      "011110101000010001000100010000",
      "010110010110101111100101011010",
      "011100010000101010100111010001",
      "111100111111100100001111101101",
      "011111000011010110010111001101",
      "001000111000000010100000010100",
      "010000000010110001110011110010",
      "110011000100000110011000111110",
      "000100110000101011000011111100",
      "101001001100010010010001100010",
      "101101000100011000110011111101",
      "110001100101101101000011100101",
      "010001001011100001111111100000",
      "101111101110101011110001010111",
      "110101000001100100001011011011",
      "000000111101011011111111000101",
      "101111111000100010100011110101",
      "011101110100101000010111101101",
      "000110111110101100111011111101",
      "010011000111000010101000111011",
      "001110011001111011100100100101",
      "011110001011011011110110110011",
      "010100010101001110101010111100",
      "000010011100000111000111000010",
      "111011001011011010101001111000",
      "111110011000011010001101011001",
      "101000100100111010101010010100",
      "111101101100000101111101100110",
      "001111000111111001010010000001",
      "001111010111000000010100001100",
      "000011011000101111100110110101",
      "100101001100000000110010010000",
      "110110001100000110010001100111",
      "000010110000101011110110010000",
      "110111000000111111001100101000",
      "111011011101000000011101011101",
      "111111110000001111100100110010",
      "011011001010100100100110110110",
      "101111001110011111111010000101",
      "100011000100001000100111010000",
      "101100111000101111110000111110",
      "111000000100101111111010111101",
      "100111111011010000000001000111",
      "110010010101010001000101110010",
      "101101101100011000001110111111",
      "011100111100001110101000001111",
      "101111000000001111001101001000",
      "110101100101101000010110000101",
      "110100011000000010001111000100",
      "101001110000110101011010000110",
      "011000110010001101110010101010",
      "010101011001010110110001010110",
      "101110111111101100010011010101",
      "011100001111010011100011101000",
      "001111110011011000010000001000",
      "001101010000011100010101111101",
      "010011111000110010111101010110",
      "110101100001011100101000011100",
      "100000010001000011000101011101",
      "001110001010111011010001010001",
      "101011111001010111100111111110",
      "111111010011111100110010000101",
      "010101110011000000000111101111",
      "101101000011101010110111010000",
      "001100001001000110101100011101",
      "001111100110011000011100110100",
      "100101110110010000011000011000",
      "011110110101111000000010110100",
      "110001100001100100100111100100",
      "011011101100101001010110000101",
      "100011001010010101101110001101",
      "001001011111001110011011100010",
      "111100101001001010010100011000",
      "000001100001110001000111011100",
      "000011100100111100011000001011",
      "001110001111101101010000110110",
      "101011010110110111000100000110",
      "000100101111101101110001101100",
      "000101011110111000011101000101",
      "010111101110001100011000001110",
      "110101111000110101101100011000",
      "011000110001011110111101000111",
      "001111000000011111010010100100",
      "001000011011000111011110110011",
      "111100110001011101000010100110",
      "010000001111000011001000001101",
      "010000100111110001000111011000",
      "001100101110001110011011010010",
      "111101000100110010011010010100",
      "001111001001100011001001101111",
      "011100111010111000110001111010",
      "110001100000101101000111001111",
      "000000011111111011100111000000",
      "000110000111101101000100110101",
      "010100011100001011010111101110",
      "101110100010010100010011110111",
      "010001111110010000010010100110",
      "001101111011100100101111110011",
      "011100111000000001010111001100",
      "101111100001011001101110011000",
      "101000011011001000011110101010",
      "101001011111000101101011110010",
      "001010101110100100011100011010",
      "111101101010000010101010100101",
      "010110110110100001010010001100",
      "001011111100011101101111000000",
      "000000011010101011101011101000",
      "110111010001101100010101101111",
      "010110101111101001101010101001",
      "010001111011111100101101101111",
      "100000011001011001110001110110",
      "100000011101100111100111010101",
      "001111001100101010010110010011",
      "011010100000011000100010010001",
      "101100010100111110100110000101",
      "100000000100001011101001110101",
      "000000010110000110110011001100",
      "101100110111101101111001001100",
      "100001111001101011110110010100",
      "100010111111110010000101000000",
      "011000011001101000100101001010",
      "101101000101011101001001100100",
      "000110100111000011101011000001",
      "100101000110011011111001001101",
      "110000000000000110011100111011",
      "110101001101010101011110101101",
      "111001111101110001011001111000",
      "000110101001010111101101111010",
      "101011011111100110001100110111",
      "001111010100110000100011001011",
      "101000101011110001101100110011",
      "111111111110000100100011011000",
      "100011001111010110100000101110",
      "100100010111000011111000100011",
      "101110111011110111000001110110",
      "001011010000001101010101100110",
      "100000010110111110111110000010",
      "100000000001010100100011000100",
      "011001101110111110001011100101",
      "010101010100110010101010101100",
      "111001101001001111101011001000",
      "010100010010000000000011110011",
      "000000000111111101010111101101",
      "110110101000100000110000001100",
      "001110000000110000110011111101",
      "111011100010100011110011100000",
      "101100110010010100101101100010",
      "111101010010100001001000110011",
      "110111100001001110000111111100",
      "001000101110000111101111111111",
      "100110011000001101100110011001",
      "110110101111110011011101001010",
      "011101000000001000111111000101",
      "110000011101001010011111001110",
      "000010100001111111101010001111",
      "110100010000101001001100000000",
      "001011110011001010111011001101",
      "101110011111111101000110011010",
      "111001110011101101010000011001",
      "000011101010011101101000011100",
      "111000000111011110011011011000",
      "001111011000110101110100111101",
      "011000000101010011110110001111",
      "111101000001010000000001000001",
      "011101101111111000101101100000",
      "010101000101001000100100110101",
      "100011110011001101001011000001",
      "111000001101000001010111000101",
      "010011011100011000011011001101",
      "111000100111100110000001011001",
      "100000101001001001100010110011",
      "001110000000010011110110011000",
      "010101111011010011101001011001",
      "100110010111101100101100100101",
      "101111010110101111000101100000",
      "110010010000000111010001010110"
    ),
    (
      "110001101001001011100010000010",
      "011100100010111000011110001010",
      "101001000110111110101010001011",
      "010011001011001010110011110011",
      "110110001000111010001011111111",
      "000011100100000001010111100011",
      "110100010001100101011111000001",
      "111110101001100110001101111111",
      "101111100000101011001000100111",
      "101110001100000111101100100001",
      "011010000011100101010010010110",
      "000011000100010010001000011011",
      "001100010100110110101101111010",
      "000011111101101101100111111011",
      "100001101111110001111010011011",
      "101010111001100110001000001110",
      "111111101110010000101011100110",
      "110000001110100010011010110000",
      "101011001000111101110101001101",
      "011001000111011110001110100011",
      "001110001001010101001100000001",
      "011010111001100110011011100011",
      "110111001000100011000101000011",
      "111010110111010011101101001000",
      "010100100110101011101010100110",
      "110110110110010110011011010100",
      "010010111001111000001010000000",
      "011000100111111111000101110101",
      "101110100101010101011000010111",
      "100011101001001011100000001111",
      "001011010000111000001111110001",
      "111100111000001111111111110010",
      "111000001010010110000011100010",
      "011001100010010111000111100101",
      "010010010011111010000011001101",
      "000001110100100111111110001111",
      "001110010011110110001000000010",
      "011110000111110010011011010011",
      "001110111011111010001010000011",
      "101011101000011110101110011111",
      "000001100111111011100101110010",
      "100111100101001101100110011100",
      "010100000010111101110010010100",
      "101110100011000100110110101000",
      "010000111100001001110110000100",
      "110110111110011110000111110110",
      "011011101000010110000011001000",
      "010001001001101000110110101111",
      "010001110110010000010000011101",
      "001110111001110010101010101100",
      "011011101111010100010101010110",
      "011101000100001111111111100111",
      "001100001111100010010111001011",
      "001000100101000101111110100010",
      "101110101010101100110010001001",
      "000111000011110000101000001111",
      "110000111110000010110101010001",
      "111000001101111001011110011110",
      "000010100000111111000111011001",
      "011001000111011001001000111100",
      "111111101111110110111101111001",
      "111001110001110110110101001111",
      "000111001110000010011001011100",
      "010100100011010101100011110101",
      "110010111111111110011011000011",
      "010101110110010101010011000110",
      "010010010110100001000011101101",
      "000011101101100110101100001101",
      "001001110000001001001011011011",
      "111001001001001110011011111000",
      "010011000111101101011101101110",
      "000001110000101010101101110100",
      "010100100010000101110101100000",
      "000000001010101111100110100101",
      "010011100111001000110000001011",
      "110110100011011010011011011000",
      "000110110101010110011010111010",
      "100111011110010111110111111010",
      "011000100001011011000011101011",
      "010100010100101010101101000000",
      "100110010111101110101111011001",
      "000001110110010010110100111111",
      "000111100111010001111110110100",
      "100100011000001000110110111101",
      "000110111010101010111000000110",
      "101001011101100110001011011001",
      "100011100010000000010010110110",
      "111000001010001110011110000001",
      "111001111100110100101101100110",
      "011011000001011100001000000001",
      "011101001100011101101011011001",
      "101000110001011010101010010000",
      "011010011001100110101111000100",
      "100001101011110001001010101001",
      "101000100111110100011011100000",
      "011111001100101011011100011110",
      "101010111010011010011101111101",
      "100100011001111111111001001001",
      "101101101100010000110111011000",
      "111001100011100111101100111110",
      "111100100101011000011000011111",
      "100000100000011100011010000111",
      "011010110011011110001000101011",
      "001110010011100110110000011010",
      "101001111100111000000110001111",
      "010000011101011101000000011101",
      "101110011111100100100000001110",
      "101110110000011000000010010010",
      "111100110000111100111011011101",
      "001100010110010000101000101011",
      "000010100001101100110010011101",
      "010110100110111000001110011001",
      "101111111110111001000010101100",
      "111101010011111101010111000000",
      "001100101111100101011001101001",
      "111001010111101011100111011000",
      "000000011100001111001111100001",
      "010010100110000000110111110010",
      "000111010001011110111110101110",
      "111010011000011000001011000111",
      "011011001101001011011110111010",
      "011001101110110000110010010011",
      "110110100010011011000011100100",
      "001001100101001011011101110101",
      "001011111011001100100001010011",
      "001100000100010000001101000110",
      "011001001110111011111100111011",
      "000011000001101001000101111110",
      "011111100110011101101100101010",
      "100101111111100101010001110000",
      "010011001110001111110100000001",
      "011100101101000100101011100000",
      "111001110111000001011001010111",
      "111111001010101010110010110111",
      "001010010011010000001110100101",
      "001100000001111101101000111100",
      "111000111110110011000111001110",
      "000010000110011001011000010110",
      "000110011111001000000001111110",
      "101011111010000001010110110001",
      "111000100000011000010100111100",
      "101010110000100010101000010101",
      "010100100101000000111011100010",
      "011000001011011100011000011101",
      "010101000110110101010001101111",
      "000111100011011111110000000111",
      "110110111110010001110110110000",
      "011101011101110010101010100110",
      "111000011001000000011000111101",
      "010110000001011001001101111001",
      "101100101111001100111110010000",
      "010101000111000111010000110000",
      "111000000010000011001010001101",
      "001010100011011101001011100010",
      "100011010101101011101001011000",
      "110101100010010100000010101011",
      "011100110011000011111100111001",
      "001111101100110111000000011001",
      "111010010111110010011011110100",
      "001110100001110011101100001101",
      "100000100001011101101111010101",
      "001011001010111101010011110011",
      "010111100101000000101001101111",
      "101100110000000001010110110011",
      "111010010100001001101100011111",
      "000101010111011100001000011001",
      "010111011010010111000111101011",
      "010000000010100011100111100100",
      "011111110001101000010110011000",
      "110011111000000100010011110000",
      "111001101111001100001011110010",
      "001100101011100111111011010111",
      "001001001110100000100100010100",
      "111100101101110100000011011010",
      "000101111011100110000010100000",
      "001101011010000111110001010111",
      "001110010000101110000100111110",
      "111111011011000001101101001111",
      "001010001011100010100100000111",
      "000000011011000100100010110011",
      "001011100111011000011011100100",
      "100011101101010110010101101001",
      "001100101001010111110011010111",
      "110111110000010111000000100000",
      "001101001111110100111111010110",
      "100011010100010000010111010000",
      "111100001111011000111110001110",
      "111101100111101110101100101110",
      "110010100001011011010010111110",
      "011110110000001001011000101011",
      "001111000100111010101000111001",
      "001101111101011111011011000100",
      "100111110110011011010011010000",
      "000100001000101000101110011101",
      "000110100111110001100000010111",
      "110000011111110100001010010010",
      "011110111011001010010000010110",
      "100101010000110001100100010010",
      "110011111111101110111011010111",
      "010100110101011110001010111100",
      "111000011010010110101001010011",
      "110011100111000000010110100111",
      "101001111110100110001111011001",
      "101110001111100011000010011111",
      "000001110111110111001111010001",
      "010110101111000100011100111100",
      "000110001000011110000011100111",
      "111010100100011111011111011110",
      "111100100010100111000000000001",
      "011101001101011010010110010011",
      "010010011011101011110000001000",
      "000000110000001100100010111110",
      "011010000100000110110111011011",
      "110011010101000010000111000011",
      "110000110001000101011101000110",
      "010000101100000100111010100100",
      "010110100100011010010110011110",
      "100000111111110000001010111010",
      "100010000101001101101111110101",
      "100110001111100111001110010000",
      "011000000001110010010000101100",
      "000111011000010101111100001100",
      "000000001011001100100010010011",
      "000101001011100111100110000011",
      "010011011001011111111111110111",
      "101001011011000110011010010110"
    ),
    (
      "001001111100010111111101101011",
      "000111010111000110011000111000",
      "100011111001010001010111001111",
      "010100000111111001010000001111",
      "010000000111101001010101000010",
      "100000001111011010000010110001",
      "011010011111001100011001011110",
      "011111000100011001001111110000",
      "101010000110101100000101110100",
      "001111110000001001100110110100",
      "000001110100100110100000111100",
      "100110110010000001010000111001",
      "001101010100001110100100011000",
      "000011110110101011001111101010",
      "010111100010111011000100101001",
      "110001011101100111101111011000",
      "101011010111011100000010111110",
      "001100100101101111110111010111",
      "110101101101100101111000100101",
      "101100111011001110000100101001",
      "000000011110011100110010000101",
      "111010010011010010110011011111",
      "000010111111001001111011010100",
      "100001001001011000111010100001",
      "100100001010001011000110101111",
      "111100010011000101010111001010",
      "110000010100101110000111101011",
      "001110011001011101111111000100",
      "101110110000101011111010000011",
      "100010010010001110100111101111",
      "101100100111001100101100001011",
      "100011100010011111011010110000",
      "001110000100100101101110101101",
      "010110000110010101000110110111",
      "000101111000100011100010001000",
      "100011000100100101000010100010",
      "100100001100111111101000110101",
      "010010110000010110000011100100",
      "101101101101111011110000000011",
      "000011101101101100010101110000",
      "101011111010111111100000001110",
      "111110100000000100111000010111",
      "010110001011010110110011000101",
      "100110101101100010100001001001",
      "010011111101111010010011111011",
      "101001011101100100111000000101",
      "101111100000101011000000111111",
      "000001010110010100010100001001",
      "010011010000111110100000001010",
      "101001001100111110000101010010",
      "001001000101001111011101011010",
      "100101001111110100011101101001",
      "100011100111101100001110110111",
      "110011111111110101011100110011",
      "000001011111001101101101111011",
      "010011101011010100101100000101",
      "010110110001000110001010010100",
      "101001110001110110001010100010",
      "010111100110011011001000010011",
      "101111010111001010001110100101",
      "011000001100010110111010000100",
      "100101011001011110000011010110",
      "110111000111111111001111101111",
      "000011001010000111110111111000",
      "100011100100110110001000010110",
      "100101011101001110000010100100",
      "011000010110111101111000010100",
      "001111110011100110011001111000",
      "001111001100010110101010001101",
      "010000001000100111011000011000",
      "010101010001111111010100101111",
      "100110111100110011111010100000",
      "101111100000010010000100101011",
      "111100000110010011100111001110",
      "101011110001000111000001101011",
      "000001011101110100000101010101",
      "111110011100100111010010100100",
      "001010111100000001111011100001",
      "100111010110110001110110000110",
      "001110101011001011011010011010",
      "100000011100001010011011000110",
      "000101101110011011000111101100",
      "001011000011011110111011010110",
      "010010101101010101011010101110",
      "011001011011001010111101000100",
      "100001010100011100100110110011",
      "101011011111001101110010010001",
      "100001010110010101011100010110",
      "010111001011110011101001010100",
      "000010101001011101001111110101",
      "101110000010100111111001001111",
      "101010011101100110100100111100",
      "111101010010101001100100010001",
      "000011110111110111110111111000",
      "110101000001100110111110110110",
      "011100110110001000111010000100",
      "110100010101000101011001011011",
      "011101111110001010110011000110",
      "000111011111000100110010001101",
      "111101001101001111000111001100",
      "100110110011100100001110001000",
      "001001011111110100000001000100",
      "000110010110101001101100110011",
      "110110010100101000100100001101",
      "111100010010011000101111100111",
      "011100101011010010000010000011",
      "010100001010000010110100001110",
      "010111001001000000100110100111",
      "100011001111100100100010001110",
      "000001110000111101011110001101",
      "101110001100001010001111101111",
      "011111001100000100100011010010",
      "111100101111101100110010111011",
      "001100011101010010000101101011",
      "111011110000010001000000100110",
      "110111101101101101000111001000",
      "110101100101001101110110100110",
      "101001000111000110001101111010",
      "000100111011000010111111100100",
      "111111010111100110100110111001",
      "000101100010111100001011100010",
      "101000110101001011010000010100",
      "111011111100011000100011001100",
      "100101001000100101100110000111",
      "011100001001110111111100111101",
      "110101001010110100101001000101",
      "000110010110101111111100011100",
      "100010010100101110100011111001",
      "010111000100011110000111100100",
      "101010011110111111001100110100",
      "100001111010011110110100110110",
      "001111010011011111010100111111",
      "101101100111111010100110000000",
      "100011110100000001001110010111",
      "011101101010110000101111001001",
      "000101110001101010111110111101",
      "110110011101011111100110001110",
      "011100101000011010000011000101",
      "110100000000010001110001010010",
      "111101110101001001000001011101",
      "100100000111110101111011001010",
      "001011100101001100010000000010",
      "100101010101111000000001011000",
      "010110101100001100110001101000",
      "110001111101010111111100001000",
      "110010111011001011011101010001",
      "010010000110100101010101110100",
      "111010010011001110000000001100",
      "110011001011000110100111110010",
      "010010111100001100110110001110",
      "101011101011001000000000111011",
      "101000101100111011111001101111",
      "000001100101000001011100101100",
      "011010001000001011001100100011",
      "100011110000111100011110011111",
      "101010101110110111110010101110",
      "100111101100100111110010101101",
      "000000001101010111111010000010",
      "000011010001110001001101011011",
      "011111101111100010010001110110",
      "000000111110111101000010111100",
      "011001001111100011100111010011",
      "110000111100011110011001001100",
      "001000111100111111110110010111",
      "001000010111101110000000011111",
      "111110100000001100010100010101",
      "001110110100111000100101011111",
      "100000001100110010111000011001",
      "110100001111000101100000000001",
      "010010110001111101010111010001",
      "100000111111110000100011011011",
      "100011101100000101001111011001",
      "111110010110100100100100111000",
      "111111111110111110010011101111",
      "111110101001111110001000100110",
      "100111100010011010011011110000",
      "100101101110110000111000111001",
      "101110111110100110100101010011",
      "111000000001001010110111101110",
      "001100111111011000010101011000",
      "011101000111100011100011001100",
      "100110101110110110101001000010",
      "111111111100111101100101111001",
      "000001000101000110010011100111",
      "100000000101110000111101111100",
      "001010100101000010111110001111",
      "100110110000000111000111000100",
      "000001010101111000100111101011",
      "110011010011110000110011101110",
      "101110001010101000111110100000",
      "011110001111100100001001010011",
      "100100111111111010111101110100",
      "110001000101110101101101000100",
      "110111111011101010111101110100",
      "110000101000010000001111100101",
      "010011001110110000101000010111",
      "111011100100110100111110001111",
      "110010000011111110100101000001",
      "101100111110101100001101010100",
      "100000110110001110110000000001",
      "110000011001010000001100000111",
      "111000010000100010010000001110",
      "111001110001000101101001101011",
      "000101110100111010001011100101",
      "100010110010111010100001110111",
      "010001111100011100110001100110",
      "111000111101100010011011110001",
      "001001011000010001111111001000",
      "001110011101010011110000100101",
      "111000011100111001111011011111",
      "100001000100001010011101110000",
      "010101110000111011101101101111",
      "000000101110111001011111100011",
      "011000101010101100110111111110",
      "000100011001001010010010111011",
      "001010101000001001000010000001",
      "111000011110000000110001000110",
      "000000100101100010110100111100",
      "110011100000001010101100010001",
      "101011100100110100111101000110",
      "101110110001111000001011111010",
      "010101110111010110101110100000",
      "000001001010000001010101000101",
      "011010000101011001101011001001",
      "111111110000001100101110110100",
      "100000010000111000011010111001"
    ),
    (
      "111111111011011100101000010111",
      "000100001110100011110011100110",
      "110011000111100101011010011110",
      "001110001111001111001010110111",
      "110001010011000011000000110011",
      "110111000100001100010111110100",
      "101100111001111111001110111101",
      "001111010101100111000111101111",
      "101110000001010110000101011101",
      "111010010011000001111001000110",
      "101101100101001111101010001111",
      "000101101101001111101001111000",
      "100110110000101001011000110011",
      "011111010011101011111010101100",
      "100100010111100101011010110011",
      "111110010110001110110101000111",
      "001111010011001101110111001000",
      "010001001011101000111111011000",
      "111101000110000011010000101111",
      "110000010100010010100010010001",
      "111010100101100011111111110010",
      "001101111001000100010010001110",
      "111111111101101100000001011111",
      "000011010011101101010100101010",
      "110100011010011111101011101100",
      "010110110010010111110100001000",
      "001111000011101010111001110101",
      "110111100101110101101110011110",
      "001111111001001110011110111111",
      "101010110000110011001000000101",
      "110101111101100010101011010010",
      "111000111001111000101101001000",
      "010101101110110000110010011001",
      "100100001000000101001111010110",
      "101100100011111000111011110110",
      "011010010000010110111000010000",
      "000011001101110100000101011010",
      "010101110110001001010100011100",
      "100000111111010101010110100111",
      "110101010110100110000101100000",
      "010000110110001101100000000011",
      "010011011001011000101011100110",
      "011011001010001000001111011111",
      "110110011101110111101100110011",
      "101011000001110101111111000100",
      "000110101100011111010010011110",
      "100111110100101011000001011101",
      "100101110000010101111011111000",
      "100110101101010100101101011011",
      "111000100000101110000000100100",
      "001110100001110000010010010010",
      "110100110000001000101011100110",
      "011001000111001101110101001111",
      "101000101110011010111101001011",
      "100101101101010001111110100011",
      "010111110100000101111011000101",
      "101011001101111001111011100000",
      "111101110100000101100001101001",
      "000011101110010001011000110100",
      "001011001100010110110111101110",
      "110000010100000010100111100110",
      "000110001110111000011111100011",
      "000010000101100100001110001111",
      "001111110001100000001100011010",
      "101000010011001110101011111011",
      "011101011110100001100001100000",
      "001011011110111101101111100000",
      "011010011101010100001000000010",
      "111110100000101001011000111000",
      "101010010101010000000100000111",
      "000010011010110010010010110111",
      "101111010000101010000111001001",
      "010111000010000000001000101111",
      "011101010000001110001000111000",
      "111111010110110001011101101111",
      "000001100100011110110110110110",
      "011001111111001010100111011111",
      "111101101000000110111001000011",
      "011100100010010010110001011101",
      "010011011000101100110111101100",
      "100000000100000101001001000111",
      "000001001110110101011101101111",
      "101000110100110010011101101111",
      "110001101011101000000100000101",
      "010111101111111100101110101110",
      "001001011000110000101111000000",
      "001111000110100100010001001001",
      "011110010000110000000110011011",
      "010111011110111000010111010011",
      "000110011101101111011011001010",
      "111010000011001111010100010010",
      "110101100111010001001110000001",
      "011011101010001011111011110000",
      "011111110011011100110010101011",
      "110101000000100000011101001001",
      "111001010001100111001011000000",
      "111000001001101010010110110011",
      "001000110001001010101011101101",
      "101011110001001111111010101111",
      "101110010010011111100101000010",
      "011001101000010011110110100111",
      "111101111001110101101111100000",
      "111100110100010101100001011101",
      "011001010000100010011010110110",
      "101001001011001100000010011100",
      "001101111111000110100011001000",
      "001011011101100111000101010000",
      "111101001001110110000000001100",
      "001100010100011001110100011100",
      "001100010101100010101010000010",
      "011001100111101111001100100011",
      "100100110011110101011111110110",
      "110111001001100001100101011101",
      "100011100011001000001000110000",
      "110110111100011101111110001001",
      "011001010010000000001111010010",
      "111001100111001011010110111000",
      "101101011000010100101001010010",
      "110000100000011101010000100010",
      "000010111011100000001110000101",
      "111001111000010100100010011010",
      "001010001111111010000101001110",
      "101101111000000001101110011010",
      "010110011000011100101111101111",
      "001110011001100001000010110011",
      "100001010110011000010110100111",
      "110111000001001001001110011101",
      "010011111010011111011010000100",
      "110100100110001011001001010010",
      "100110110011011000100010000101",
      "100010110111011111011011010011",
      "110100101110001001111100000001",
      "010101110000111100011110100100",
      "111111101010100111000011101110",
      "101000111100111011100001100001",
      "011000011011001101011111110110",
      "110001001101011100001001100110",
      "110100111100110001001000011000",
      "101000110101111100100000101010",
      "101001011011100101111000010000",
      "110011110100011100111000100100",
      "000001100000000110001000101110",
      "001110100001001010110110001001",
      "011111110100101111110111011010",
      "100100100101011110010010000011",
      "001101111011111001111110110000",
      "011010101001001100100100100011",
      "100101100110010111000011101001",
      "001001011101110000011001101111",
      "011010001110011100101100010111",
      "011101110101011001100110011100",
      "001000111001101111010010100111",
      "101100111000011001111110100100",
      "011111011001110101011101111011",
      "001100100111111010100001001101",
      "100000010110101100111011101001",
      "010110001111101100100001111110",
      "101011100010101100011111000111",
      "001100101001001010111100001001",
      "010110101010100111011011001111",
      "001010011001101000101011010110",
      "100010111100111110110110100010",
      "001100011000100000111101111101",
      "110100101010000111101111011100",
      "011101000011001110101000011001",
      "010110100011000010000000011001",
      "001011110011100010011110011001",
      "000001011100010000111110100111",
      "100011101111110111101010100000",
      "010101010111110111100111001110",
      "001010111000101100100000110001",
      "010011111100101001100011110100",
      "111110111000001010111100000101",
      "010001001111111100101000100010",
      "001000100000111011011010100011",
      "010101111110000010000000011010",
      "100100100011010010111010010100",
      "010111101001011000100101110110",
      "101111110100110111001000001101",
      "101010101011001110100011110111",
      "000011011000010011011101010011",
      "000111010010101100000001000001",
      "010011010011111001011100100111",
      "111111010001010000111001101100",
      "111000110110000101100101001001",
      "100110111010001110011101101111",
      "001100010110110000011111010111",
      "111010010011000100111010001100",
      "000011101100010011100000011011",
      "100011100010110011111100110000",
      "101011011011011001110011100010",
      "001000001111100001110001101111",
      "111101101100011101110110010110",
      "101101110011001001010111110001",
      "001110110011101110101111110010",
      "001110100001000000111000100110",
      "011010101000000110000010101010",
      "111101111101110111111010100001",
      "000110010100100100101111111100",
      "000111110011010110111010000001",
      "101101001100011110000010011101",
      "111000000110001101001010000111",
      "010010111011101100111000001010",
      "101100110101111110010000110110",
      "100110011010101110100100011111",
      "111010010011110100101100000100",
      "011111111110001001010001001110",
      "100111011000011001000010101000",
      "010100010101000001000100110111",
      "100110111001100110111100111001",
      "011011101010001010111010110010",
      "100100110000000001110100000111",
      "100001011101001000000010001010",
      "011000000001101011000010010011",
      "010110001001100000001001010110",
      "010111100011011100011101110111",
      "000001001000110010000000011101",
      "000111101101100110100010101100",
      "100101101001100000001001001111",
      "011001001110110111001010011100",
      "111101000110101000110100111010",
      "000100000101001101110100010001",
      "001001010000011101000010110010",
      "001000001110111000101101100000",
      "000010110111000010110010111001",
      "010101000100110110001010000000"
    ),
    (
      "110111100000000100010011001000",
      "111100000011101101011100001111",
      "110101110100000100010110010111",
      "111111110101010101111001100000",
      "000111100010100011000010001001",
      "011001100111010101011001010000",
      "010101010001000001110001000010",
      "011000010011110000101110000100",
      "111010101110110001100100011110",
      "001001100110001000110000011001",
      "011011100001111101001101011001",
      "110001010001101010111110100001",
      "000010110001111010100101110000",
      "111001100110010101111101010011",
      "010011010101001111111001000111",
      "100001100110100011101111011011",
      "100111110011010111001010001011",
      "001010011011000001001001100100",
      "000101101101110111110100111110",
      "001100110100111010011011100100",
      "101111001010111010100110111010",
      "111000001001100100110011111001",
      "101011010000100110101010100111",
      "111110100000100101000010100011",
      "000111010010001000011101001001",
      "001101101101110010100100011100",
      "110100100011001011000011001110",
      "001010111010100010010000010010",
      "101000000111011010001000001110",
      "110001100011000110001101100010",
      "011010101011100001010010000001",
      "010111110100100111100110100111",
      "010001001111010010101100101110",
      "101011011001001010110001001101",
      "110000101111110011101100111000",
      "100110010001100001110011100001",
      "100010000001000001000101000000",
      "101000110110001101100101110011",
      "011001100010001000001111011000",
      "100110101110111111000001111110",
      "101011101110111011101001101100",
      "000111000010011100010011011011",
      "001000111010111011110010011100",
      "001000001011000101101010110011",
      "100001111110110001000001110110",
      "110010010101100111101100000111",
      "001100000000011000011110111000",
      "111000011101000011001011011101",
      "100111101101011111001011001011",
      "101011000001101101011001010010",
      "101000010000110000111101100111",
      "011010110100110100011100010100",
      "110111100001010011101011001111",
      "010010111010111101010011101011",
      "000100001011100111010101111001",
      "011101101110111101011011001110",
      "100100100100010010011100111010",
      "100100101110011110011101111100",
      "100011111110000110001100101010",
      "100010101111111011000011000101",
      "010110101001110001100010000000",
      "010100011010001110111111100001",
      "010001000111110010111011001101",
      "101111100101000010011000001101",
      "110101111111111110011011000111",
      "000010001101010010001100010010",
      "011111101010010000011000011100",
      "110001000000001110111001111101",
      "001110111001100111101001110100",
      "100001110011100001110111110010",
      "011001001111101110101010110001",
      "011000101000010000101111001111",
      "101100101100101111100000011111",
      "011011001111011100110010101011",
      "100110100011011100100010000101",
      "100101010011111101000001100011",
      "111001111100001100110101001110",
      "010001110000110111101101000000",
      "010101111000001100010001111101",
      "101101101101111010100110111000",
      "110000100000100110111101110010",
      "110010000101111011010100111001",
      "011001001100110100010110011001",
      "100110111001100100001111011110",
      "111101110000111100111100000001",
      "101000100101011111011011011011",
      "111110011010010100110100010101",
      "011001011010100101000011101100",
      "111110101001100100110001110011",
      "010000011110111100110101101101",
      "000101111001000110011001110100",
      "101111011000100011001011000110",
      "001101011110001111111001110100",
      "000111010101100010111111000110",
      "001010110111110110000000110010",
      "101000011110100110111000011010",
      "100100011110011110101010010100",
      "000001001110010111111011110101",
      "010010111000110011011001010010",
      "011101001000010100111101111101",
      "110010111001011011000001010010",
      "010000111001000010000111111011",
      "101110000001000011110011010101",
      "100100101100001111110000010101",
      "100001001110111111110100110100",
      "010101101101010001101001101001",
      "100111101100001010100010001110",
      "100011101010010011111000000010",
      "101101111110110010110101010001",
      "001000111000111110011100011010",
      "110100011111001000010010001010",
      "100101110101001011110100111110",
      "101101101000101101001011111100",
      "010010110101101001000001010000",
      "001001110011000110101010100000",
      "101000010011101111010101001010",
      "011110110001001011010111001000",
      "111111001010110100000101110000",
      "000011010111010111100000111001",
      "010001111101010000101110011110",
      "001010101101011100101010010100",
      "001011100111111001101100100110",
      "100101110011100000011010001100",
      "000001011111000111010111111000",
      "100100101110110111010101000100",
      "101101111101101000101101110111",
      "010111011101101110110100101000",
      "100110000111001110010001100110",
      "110111110010110000000011001110",
      "000011010000011101011011110001",
      "011011101001000011000111010011",
      "010000000000100100111001110110",
      "010100101010100000110001001011",
      "101001011011000101010110111110",
      "101000101100110110010010001100",
      "000000000110101000100000001010",
      "111011011100100010001011111101",
      "101000101101100011000001100111",
      "001101001110011000110001111111",
      "000100100101110110011010101001",
      "101110000110001100001000000111",
      "100010000111110010110100010110",
      "001010111110100001011101000101",
      "111111011100001000011010011001",
      "110011000101101010011110000000",
      "010001010101010001000011000101",
      "110001111100011111101111011001",
      "010000101001100000100000100001",
      "111010001100000100110101111101",
      "110100100011000011100101001101",
      "001111010111101111010001001001",
      "101000000001010100001011110010",
      "000001000101100100001011000111",
      "001100101000110010110000000000",
      "110111101000101010011010011010",
      "010011111110011010111010101110",
      "011101101000110010010000100010",
      "110110010111110000100000101001",
      "000011000110101111000111101111",
      "110110110000100010110011110001",
      "111010101111111010011010111010",
      "101000011110011101001000000010",
      "110101000011100110001010110101",
      "011111010010011110000000000101",
      "100100100100000001001100000011",
      "110100111010010101001101100100",
      "101101001000010000010110001101",
      "000101111100111010001011100110",
      "011101101000000011100011100010",
      "111100100100101000100110010000",
      "010011110110000110110001000100",
      "001101101101111111111011110101",
      "111011000001101011000010010100",
      "011101111110111110011001001001",
      "011101001001010011010000110011",
      "010001001100110100011110011111",
      "000111101110000011110010000111",
      "001011001110110110101001010110",
      "011001010000001001010111001011",
      "111000111001001101001001100101",
      "100101111111011000101011001100",
      "000010110111000010100000010101",
      "000101010001001010110101100010",
      "100000000101010000101111010000",
      "111000010011111011111000101100",
      "000101010001110101001111000001",
      "101000010010111110100000101100",
      "010010001000001000001100111101",
      "001101101100111111111110011101",
      "010101010110111110100000010000",
      "100001101011001010101111110010",
      "110101100001111011110111111000",
      "101110111100011000001101000101",
      "001110100110001110000111000100",
      "001011000111100001001110001000",
      "110111010101011000100010101001",
      "010111100110110110001000101001",
      "101010000111100111000011010011",
      "000110000010000001001000010100",
      "110101000100001001010011010101",
      "011110100101000101110000101000",
      "101001001100010001110111101111",
      "000011010111010000110110011101",
      "100110011101001001000000110110",
      "100000010001000010100101000001",
      "101010000111000100100010010111",
      "110011010010011010100000100101",
      "111010010000111110110000010110",
      "100011001110000110000011111110",
      "000011011000101001110111011001",
      "100100000010111010001011101110",
      "010101101100001100001010101111",
      "000101001001100001111101100100",
      "000111010010000011001100011111",
      "111100001101011001101111001110",
      "010001010001000101101000010110",
      "001100111001000011011110001111",
      "011111110100100101011100010110",
      "111111010101101111100001000101",
      "010101000111111010010000101110",
      "110001110110001100111011001000",
      "110011010011110111001111010011",
      "011010100001011010111001000100",
      "000010000000010111101101111110",
      "110100110101110001001010011000",
      "101010110111010001111100101010"
    ),
    (
      "100010110011001011000011010010",
      "100010000101000100000110100110",
      "011010110110101101000110001110",
      "110100000010000010001101101101",
      "010010111001101111000000100010",
      "010011100111111000110101000000",
      "110110010001010111010010010100",
      "110101101010010000011110001101",
      "101101011001110010101000010001",
      "000011001100101000111001110100",
      "000111100011110001110100110110",
      "101001111100111001110010010011",
      "010001001000100111011110111001",
      "100000010011111111000101100000",
      "111111100100111011000000000011",
      "001010000011101110000100101101",
      "100011111011010111100101011101",
      "111011010110000000001010100100",
      "011101001101011100000011101000",
      "111101010011110111011001000000",
      "001110111111110001111111010100",
      "000011011110111011001101110101",
      "011000101111000111110111100001",
      "100000111011001001001010101110",
      "011110001010100010110010011000",
      "000100100110010001110001000001",
      "110100111001110011100111001110",
      "100110101101110010010101110110",
      "110110010100110010010100011101",
      "000100011010001110011010111111",
      "100010010110001001011011101000",
      "000000111011001101001101111100",
      "111011101110111100000100011001",
      "110011110110000101100111101001",
      "110100001001111011000000111110",
      "110001111100000100000011010111",
      "001110010001001111000101111001",
      "010010101000111100011001111101",
      "100011110110000001001100010101",
      "001011010010101011001100111111",
      "100001010000111000101001010100",
      "111100110100010001111011100010",
      "101111011001000010010100011110",
      "111010001010010110001100111101",
      "110000011010111110110000010101",
      "000101011110100111100001011001",
      "101111010100100010111001110001",
      "100011011110110110100110000010",
      "110011000110010100000010101101",
      "101000100011110011000010110111",
      "000010111010000000001111110101",
      "111100101010001111100100001100",
      "011000001001110100100111100110",
      "011000001110111101000001111110",
      "000101110010110010101111011100",
      "001000110101100110110111100110",
      "111001011111010000101000010001",
      "001101000110110111010100100000",
      "000001001010001000111011011000",
      "110110111001111101010111010000",
      "110010100111010110100010010101",
      "101011001000010110111100100000",
      "100111001111000101101101110110",
      "101011001010000001001010100010",
      "011000011100100001001111101101",
      "101001110111010011011101010101",
      "001001000100110110011100011011",
      "100000111110011101001001101100",
      "000101001101101000111100100111",
      "101010001001001110010100000001",
      "001001101010111010011111010101",
      "111001001100110100110001010011",
      "111111011111111101011110001111",
      "010111011110111111000011101101",
      "101011001110000101011111010100",
      "010010000001111001111100010000",
      "101000110010110011111100100000",
      "011010001100100111010000110010",
      "010100110111011000000001111011",
      "100011101111111000101011100001",
      "110101110001100101101011000100",
      "111001000111000001110011101000",
      "110011010000100001110010110011",
      "100000101000010000011110000000",
      "110100111010110111100101001100",
      "010010011101111100100111010001",
      "100110111110111011101101000010",
      "010111000011000011000110011001",
      "111111000111011111000000110100",
      "000001010110000001101000100100",
      "110110110110100100111111001110",
      "111101111111111010001111011101",
      "011011010100110100000110110101",
      "000111100110010010010010101010",
      "011100000100111011001000101000",
      "011010111100111111010100010001",
      "001111010001100111011110111110",
      "101000110110011010011110000011",
      "111010110101110101111111000011",
      "000000111111010101111010110100",
      "100000100000010001110101110001",
      "011001011000010111001100110011",
      "110110110011011100110000101101",
      "001010110011111000100001110001",
      "001100011101111110100111000000",
      "011111110010110011100100101010",
      "111100111010111001110011101110",
      "111001100011001011010111101110",
      "100101101010100001010111011010",
      "001001011111101100100110001101",
      "100111001110010101000101100010",
      "010011011000101000100111101010",
      "010011110000111111011010011110",
      "000010111100111100111100010001",
      "101010010010000100000011100111",
      "010011101001101101111110010011",
      "011001010101111101101100010011",
      "110000111011111101011110100101",
      "001111011101000110110100011000",
      "001010001001000101001010010100",
      "010110111001110100000101010100",
      "101010000111000100011010001100",
      "101000010101100010110011010011",
      "100110100010010010011001011000",
      "111001001100111101000011010110",
      "111000100100100111100010010001",
      "111000000101010011001100000110",
      "110111000000100001101001000100",
      "011100111010101110110111000101",
      "010001000011110000110111010110",
      "101000111001001000000011100110",
      "110000001100100000100000010100",
      "010111101010110011010101011000",
      "100111011011111000000011010101",
      "011100101101111011100100111010",
      "101000110000011110000101010010",
      "100100001010110001010110000011",
      "011110000101011011000011111111",
      "110110011110111001110011110000",
      "101100100000101011010000111000",
      "111000101001000111011011111101",
      "010011000101010100110010000111",
      "101010000100011101111010100100",
      "000011001011011010110011101111",
      "010011001100011001000110111011",
      "100011001110010111111100100110",
      "010110100010001000111100010000",
      "101111001010001100000101000010",
      "011011000001110000111001011100",
      "000000110011010001000111111100",
      "010000100111100100001001110010",
      "010110100011001100001111001101",
      "101101010010101101001001101000",
      "111100011110101011111110001000",
      "001111101100101000101110010100",
      "110010011110100000110011011101",
      "011000010101010101010110100101",
      "111001101110000001111010101100",
      "000110011011001110101100000001",
      "000001110110100100001011010101",
      "001010111101001100110011001111",
      "001101010011011100100000010110",
      "011100111001101100111000011100",
      "101101011100000111011011101110",
      "001110000111010011011001000101",
      "001100111110110111111111110001",
      "010100100011111111000010111011",
      "010101101110111000100010100110",
      "110100101011110111110100111001",
      "111111011110101101101101000100",
      "010110100101101011011100011010",
      "100000000110101001010001101000",
      "010101100101110000000111011000",
      "011101000000100100111110001100",
      "100101101001100010100011000010",
      "100110000100100111101100001001",
      "011010000001001101111011010110",
      "010111000011001011100000110110",
      "000101101101010100000100100100",
      "011010010001110011011101010000",
      "101101101110110001001011110110",
      "010001111100101011100011011111",
      "110011000110101001101001101110",
      "001010001010010011100110110011",
      "110001010110001010101110010101",
      "000110110011101011101010100110",
      "000011110101101101011000010001",
      "111100011100011110100011011001",
      "001100101010001100111000110100",
      "010011001100000110101001001001",
      "001000000111011100001010111101",
      "010110001110001101101001001001",
      "010110101001101000111101101110",
      "001000111101110110111111100001",
      "000111010000101110110111111110",
      "111101110100101111100101001100",
      "001000100110010111000100111101",
      "101100011011000111010010011101",
      "100011011101111111101100010110",
      "001100000111101011101011111110",
      "110110000010111000001001000011",
      "110111111001010011101101110111",
      "001110001111010011010111110000",
      "001010001010001111101101010100",
      "111101010100101110000110100101",
      "000000010011010111111000011100",
      "010000111011100100101010110000",
      "001010100100101100100100101110",
      "001100010101100101011110010111",
      "100010001001111011010010011010",
      "110101111101011000111010101011",
      "011111100101011001010001111001",
      "100000010011100000010001100111",
      "010010101000100110101010010111",
      "101110111101110001000000101100",
      "010100110111000101111110100110",
      "101000100001001000101110110011",
      "011110111001011111010100011100",
      "100011010000000110100101000100",
      "001110100100000111011010001011",
      "111011000000001110110010001110",
      "100000110010000010010100110011",
      "110101110001001001100000000100",
      "101101010110100001101011110001",
      "001001011010000101001010100100",
      "101011010110001001101110101100"
    ),
    (
      "010001001110011101101111011001",
      "000001101001110101111100111010",
      "100000010110100001101110100010",
      "000101000011001100000111110110",
      "111110010110101001010001000011",
      "010111011101111001001111001100",
      "110111001000011000100110010010",
      "011000010011110011111011010010",
      "000100001110010001001100111000",
      "010001010110010010110001101001",
      "110101001010010111110000101001",
      "110000110010000000111100000010",
      "010101101010101100111110011001",
      "111101000011111010110100001011",
      "011100101011110100011001101000",
      "011100100011101010111101101100",
      "001111010001001101011001110100",
      "111110010110011100101011001101",
      "000100101000111100000100100000",
      "101010011100000100010110000001",
      "011110110100100110100101111000",
      "001101101101100011000100111111",
      "100000010111110010001010010010",
      "001001010010011001101001001011",
      "101010001111110100000010111011",
      "000001110001011110011100101011",
      "000110001100011011110000010110",
      "111111101011111101100101001000",
      "100011100101001101100111000010",
      "010110010100111110111100000001",
      "101001100111100110010101110000",
      "000110001000100001001111001010",
      "111101110100110100000100010010",
      "010000110010110000011111000010",
      "000010001011110011001111001000",
      "011000011101010111110010101010",
      "010101001001010100110000000010",
      "111101000110111101001110110110",
      "110001000100100111010110100001",
      "000101111111000011111001011010",
      "100100001010100100101100111011",
      "101001101111110011010101111010",
      "011011001111110001101010001100",
      "011100001101000111001000111001",
      "001011001110010001001011110111",
      "011111001000011110111111100001",
      "001111100010101001001010100011",
      "000000010011111010110100100110",
      "110011110100110011110100000110",
      "110111000010010011010111001110",
      "100101000011100010100110000101",
      "111111110110000010100001100000",
      "110100101001011000000100110101",
      "101101111010010010110011000101",
      "011111110001000001001111101011",
      "100101011110010110110111010110",
      "100100111111001111110010111011",
      "011011000100001010001001111101",
      "100001001001110110010000100010",
      "111100100001100011110101100010",
      "010110110110110001110011101101",
      "001011001100110111111011001001",
      "110100111011000111011110110001",
      "011010000110110011011101000010",
      "100011110001000110111010101000",
      "000011001111100101101101100101",
      "010011110110111010100001011000",
      "011101010100011001111101111100",
      "000100010011101011101100100111",
      "010100011010001110100101011010",
      "001011000111110111001001001000",
      "100100011001110110101101101101",
      "001011001001001110111110111110",
      "111101100101111001000001010001",
      "100000101000110000010110101001",
      "010100110111110000010001110011",
      "000111101001010111000000100101",
      "011111111011010000000000110000",
      "001001111101000010101000100000",
      "010000010001000000110100110011",
      "011100111001010101011000100110",
      "100111100111110011001101000110",
      "100110001101011010000101111110",
      "010101010111011011000110000110",
      "110111111011000101011011100001",
      "011011111001100101010100001010",
      "000110001011111001111010111001",
      "100000111111001010100100100011",
      "010011001111010011011001111101",
      "000011010111101111000001100010",
      "011100010001111011111101100100",
      "011111010110011000000100011111",
      "001010110011100111000110001101",
      "101010111111101110010011000100",
      "100100100001011001110100010011",
      "001111100101111100000000100001",
      "000111011110001101111111111011",
      "010100001111111100000011101110",
      "101000001111110110010111011001",
      "011111101010011110010001000001",
      "000011010000011000100101110001",
      "111110001001111000100011110100",
      "100101010100100010111111100000",
      "010011100011101110011011110011",
      "010011100110011010000000011000",
      "101101100100110010011100010101",
      "111111100101100001001111110011",
      "110010100000101000101111001001",
      "111110111011010101011100111000",
      "000100110011110000011111001100",
      "010100000111110100011011100110",
      "100000000010000101010010001110",
      "110101110111110101110110100111",
      "011010011101101110110010011001",
      "100100110000110000010010111101",
      "011011110000010110000000011101",
      "001011000101010111111001110100",
      "001001100001110011001001010100",
      "000001000000001000101101110000",
      "101111111011100100100000101010",
      "000110001101111111110110001001",
      "100001011011001001101111110110",
      "101011000100010111111000111100",
      "111100011010011001000001000110",
      "010110010111101000111010011100",
      "101110001011010100110001011010",
      "001100001011110011100100000011",
      "001001101010000001010111001010",
      "011100001111101001110101111111",
      "001000000111000000011000111111",
      "100110001011010011000000010100",
      "110011100111101010010110010100",
      "011111101110100001111100101100",
      "100111101000000010100100011001",
      "001101111001000101001100111011",
      "110000010101011110010100011101",
      "000110000010010110010001001001",
      "001101111011001010000101110000",
      "010110100100111100101101000000",
      "001011000111100101111001011110",
      "100101101100111101111011000110",
      "111010110010000110100001001111",
      "001011011011010101111111010000",
      "010101010111101101000001010111",
      "011100011100010001111011001001",
      "111101110110001101110111111001",
      "111111110101000000000001110110",
      "000001101100100000000011000011",
      "010100110011111011111011100111",
      "101001111111111010100101100101",
      "111000011001010110110101010010",
      "001001100011101101011001011001",
      "011101100001011100110000100111",
      "000011111110001010000101110010",
      "000000100111110100100101011101",
      "010001001010101011011011111001",
      "111111000001100110111100000011",
      "011111011110111000101100110011",
      "100111111000110101011000101000",
      "011011010111001101001101010100",
      "000011001100101000111110100000",
      "011010010110011000101001100111",
      "011010000010011110000000100100",
      "100000001111010100111111100000",
      "010000001011111011010110011011",
      "001100101101111011010111110110",
      "100001110001010110111100010000",
      "010010010100000100011110010111",
      "011101001001010101111101101111",
      "000000001110111011110011100110",
      "011110000000010101000101101111",
      "000000110100100101111000000111",
      "111010110100000110101011101110",
      "001001000000101110111001100100",
      "010111101010010000000101101100",
      "111011110110111000011011001000",
      "111000101111100010010000100111",
      "011111000010000100110001001111",
      "011000111000010111100001010000",
      "001010100111101111000100011000",
      "011000010010010010010101011001",
      "011100111101001010111100001110",
      "000101101011000000101111000011",
      "110011011110001001101110000011",
      "001000110101100011111000010010",
      "010111011100110000111001010010",
      "100000001001100010011110111010",
      "111011010101000111011001101110",
      "011010101111000010111110010000",
      "001110001101101000111101010001",
      "110010100111010101110101110010",
      "010011101000111000000111010010",
      "100100010010010101011010101001",
      "111010000100100011001000100010",
      "110010101111011010011110100111",
      "000011010100110101100101011010",
      "000101010011100100110101010010",
      "000011000111001010001111110111",
      "101101001100100011110111000010",
      "000010101000010101000101011010",
      "101101111111000101110100110100",
      "011011110100001110001101010010",
      "100011010000001010011011110010",
      "111110111101101011001000010011",
      "010110001100111101100001010001",
      "000100010010100110001110110110",
      "110101110000110011101000110000",
      "010000010011100001110000111010",
      "001000111101111001110100110111",
      "001001010001000010011110001101",
      "011110100000101110001001110110",
      "011010010110011100001100100101",
      "010010100111111110101000111011",
      "100100000011101010000110100101",
      "011101111100111011100110101110",
      "011110000110000000010100110100",
      "011101101100110101110100011111",
      "000111111101110010010011010101",
      "111101010110101010110101111110",
      "100110000101000001101010000001",
      "011100000010110001000110011111",
      "111000000000011111011000011101",
      "111111111100101101110111110100",
      "100010101101111000010000001001",
      "100010110001100010001101100110",
      "111100110100000101010001100000"
    ),
    (
      "100001001101110011110101111000",
      "011011111111001010101011010000",
      "000111011010101101101001110101",
      "100100110101100000101000010110",
      "110100000001100100111001001011",
      "101000101100000000011111101010",
      "000100111101111111011000010011",
      "000010111000100001110100100110",
      "011010010110111001100011010011",
      "010101110011111110101111100000",
      "001010101101101111111111000010",
      "010110101000000100100000111010",
      "101110100001110110101101111000",
      "110111011001010010101010111110",
      "110010011101010100001010110011",
      "110001101010011110000011001000",
      "100110000010011011110111010011",
      "000100111000000111000111011110",
      "110101111001100000101001101110",
      "111000111000101101011000100110",
      "000010000010000111000111110101",
      "001100101000101010100111001100",
      "100110110111101100100110110000",
      "111000101001100100100101100001",
      "011011101101101111111011011000",
      "011110000011011000010100001111",
      "011001010010100101011011100101",
      "001011101111110000110110000101",
      "111110110011100111010100101001",
      "100000110111110010100011011111",
      "001101110111101111011110010000",
      "010111000111010011000110000111",
      "110010010001011011101110101100",
      "000100101100111010111111000001",
      "001010000010010111100010110100",
      "011000010100100111111010110001",
      "101011101000100111110010111010",
      "100010000101100101001000100101",
      "100000001011100001000011001100",
      "100101010101001011101000010111",
      "001001100110010100100001000100",
      "010000101000100011001000011010",
      "100001111101111000000011011111",
      "100110101101101110011110000010",
      "101101110111000110001110011111",
      "010000100001100000011100001000",
      "010111101101110011110100000000",
      "111110010110100011111001111010",
      "110110111110000010000011101101",
      "111010010111111111010111010111",
      "100101001100001011010000110010",
      "011101111000100100110100111001",
      "010110110111001000110111101010",
      "100100000011101010000010011001",
      "100100000000110101110010111011",
      "011011010010000110011111001110",
      "010101010100110011000100000010",
      "001011100101110111000101011011",
      "100010010000101001100001101000",
      "001011100110100011101010000101",
      "101100110101010010010010111100",
      "111100101000101000000001001101",
      "000010011101010111010110010010",
      "101110010000100111111011001000",
      "110011111010110100001101101000",
      "000010110011110111110010101011",
      "100110111110100100100001001010",
      "010100101000101001001010011101",
      "001001111110001000101011101010",
      "010100001100010010111110111001",
      "110000101011110100011001011110",
      "000000100000100100010001001010",
      "101110011010101000100011101010",
      "111000000000111110011000010101",
      "000101100011010000100100000010",
      "011000100011101011100001000010",
      "100011000011001100110100001000",
      "011111000000011000000010100000",
      "100010001001111010011001000000",
      "000011100111111010101100010001",
      "111101100010110110101000100010",
      "001011111100101111000111000001",
      "110101110100111101011010111011",
      "000111100111110100101010010101",
      "100010110110110100010101001010",
      "011111111011111000010001100110",
      "001111110101011111101001111001",
      "111100111101110101011110011000",
      "001001100110110000111110000001",
      "101111001001110001101110000111",
      "010100000110011100101111000001",
      "010010111101001101110100010010",
      "101111000001110100000100110100",
      "101010100000100010111010000000",
      "101111000100011111100100010110",
      "000011101101010010011111001110",
      "001001001010010001101001001110",
      "111001011110001111100110001001",
      "011100110001000110001010101010",
      "101100101111010001111110101111",
      "111100100010010001100110101011",
      "101011010100011110100111101001",
      "001100111110011110110100111001",
      "110001111010110010001000001101",
      "010100100010100000100000001110",
      "100011011100010011011100110010",
      "111101101111010100001101111010",
      "100101000000001011100100011110",
      "110101011001000011000100111011",
      "011110011001100100100000100100",
      "101010111110001000010111100110",
      "010110001010110001100011110100",
      "001101000111011101010000110001",
      "011110111001010010111111101100",
      "001001001100110001110110011110",
      "011111001011111110011000101011",
      "110111101011010011010001000011",
      "111111100111111111100110101111",
      "100110111101110110010000000011",
      "010001001000010010001000010010",
      "000010011010100111001101111001",
      "000111101111111100011010100000",
      "101011110100110011011100100010",
      "101100010111101101011101000001",
      "010110010011111010110011011001",
      "000110001010111100010010010011",
      "101111011011110110110100110111",
      "001001101010010010001111000101",
      "111110010001011101001101111100",
      "101110111111010100110100000100",
      "010000110110010010111010110111",
      "100111011011010011010001010010",
      "110111000101110111111011010111",
      "111000010011010001110000010001",
      "000000001001111110100100110100",
      "011011000010100101111101101011",
      "101100110010110101010111001010",
      "101111110110100000111010000110",
      "101110000110010100011111001001",
      "101011011111001001010110100111",
      "111101110000010101111000010111",
      "001100111011000100001111000011",
      "010011101101000000100111111001",
      "011011111110000100000000010111",
      "100111101110101010110100001011",
      "100110110000000100101110111101",
      "100101001111000100001110000100",
      "111100001110111100111011110111",
      "001011101101101111110101010010",
      "000111010100001111010100111011",
      "011101001101100110101111011110",
      "000010100010110011100111111110",
      "001011011010010110110000110100",
      "100010100000100101101000011011",
      "111100001110001101101000000101",
      "010110001010000001011101001100",
      "001101111010111001011010001000",
      "000111100101011010110001101011",
      "100111100010100111111100100000",
      "110000010010011100010101010100",
      "010000101001111001000010011110",
      "010011100110100001001111101000",
      "010111101110111001100110111111",
      "010011010001110110011011110100",
      "100111111101000011111100010011",
      "000101010000111001101000011110",
      "000101100000001111001110101000",
      "001010101100110111011110100011",
      "101001101111011001010100111010",
      "001001000101101011110111011010",
      "100000010001010110010000000101",
      "101010011000010011001010011000",
      "111001010110001110100100001100",
      "011000111110010000001011101010",
      "111001111110111011100001111101",
      "001010010111010011011111100101",
      "111010100101011001000000011000",
      "010100001111100111111110011001",
      "001111000001011011010011010100",
      "000001010111100011100110101001",
      "011111000011101011101011110000",
      "000001001100000001101010010111",
      "100011011110100010111011111010",
      "100010001010101000000001101010",
      "101110101011000001000100111101",
      "011111100000110111000000111001",
      "001111100001100100101110010011",
      "001100110000101000111100011111",
      "101111100100100111101101100110",
      "010011101101011100011111001100",
      "100100111010111101100101001111",
      "011011001011011010110010101000",
      "110101011110011111110101010101",
      "001101000110010001111100101001",
      "111101010011100110110100000010",
      "011000010100110001010111010100",
      "000010000011000101110110100111",
      "010001100000010100110110001111",
      "101000000010100011100111101100",
      "100111000001111011001011001011",
      "101001101100101011011110100101",
      "001001001001010000100111000001",
      "110101110110011010011000100000",
      "100110111111001111001101011000",
      "100001011011011001110001001010",
      "100111011111110100011000000001",
      "000010110110011011010000110101",
      "001001010010000110110011111010",
      "110001000000111001111001011111",
      "010001001000011001101011010101",
      "001110010110110011101110110001",
      "001101001011010001111000001110",
      "011110111110110000000111000001",
      "101011110000010001100100110001",
      "110100111111011110001010110100",
      "001101010010100100111000001100",
      "001101100010011101011111111011",
      "001100111000001011111001100011",
      "111101000010110111101000010110",
      "101010111011011101110101100100",
      "001000110001111110000011100001",
      "010101110110111010101101001000",
      "110001101001001010111101001111",
      "010001111101110000111001010000",
      "010101011010111101000000011100",
      "011101101101101100110111110100"
    ),
    (
      "110000011101101111010100111101",
      "101101101001000000110001010001",
      "001110000101011111000100000110",
      "111101101001010100111101011000",
      "011011000100010111101001100000",
      "011100100000001100101101111001",
      "101011100110011000000000011010",
      "110000000011100100001001001010",
      "101111011011011111110111001010",
      "010101100011010111010000000011",
      "001000010001011111100111010001",
      "101100000000110110110011110100",
      "110111111100001101010101101101",
      "011011110100000100100110000111",
      "010010011111001000011010000110",
      "111111100101110011111010001000",
      "001000101010010001011000100111",
      "000101111111101100101100101010",
      "111011010011110010000101101010",
      "001001100000011100011000111011",
      "000000101011111101001101111011",
      "001011001011011011111001111111",
      "110100010010000011110111000011",
      "000000010100000101101101100111",
      "001010111010111101101000011010",
      "111101000100101111011101001101",
      "111011110011010111100101100100",
      "101110110101110010010011010101",
      "101010100111111110010110001011",
      "001001100100000001101000010000",
      "010111100101111000001000111001",
      "111110010101001001010010001111",
      "111001110001010111101011001110",
      "011010000001111100010100110100",
      "011101010100011100101000011100",
      "011010110101000010110011101101",
      "111110100111010101111000001001",
      "110111001000111010100110001011",
      "101000111111010101100000110000",
      "010100101100101110011011000110",
      "101001110101101111101100110100",
      "100100101011001101110111111111",
      "101011101011111000100000010011",
      "100001011000011110110011110100",
      "100111110111101011000000101100",
      "000101011010111010111100010111",
      "110011011100111000010001100001",
      "001001100110011001000111100010",
      "001001110011111111010010110001",
      "010001011110111100101100110111",
      "000110010111110100100100110110",
      "011100011100011110000110001101",
      "110010011100000000110100000111",
      "001011000000101100111111000010",
      "000001011000011000111010010011",
      "110101100010100011000000010000",
      "011100110101100101001100110001",
      "010011011000111100100011111010",
      "000011111001100100111010010101",
      "010100110101110010110111001110",
      "110111010000101111000000011111",
      "111000101100101111011011100110",
      "010011000000011110001001111011",
      "001011000111100001000101110100",
      "010110010111101010011000110000",
      "100011011000001111011111101111",
      "011110111110011001010001001110",
      "110010001011011010111111010010",
      "111101010110110110010001110110",
      "000010001101011011110100110110",
      "000011110001001011111011001101",
      "101100111111001110010010000110",
      "000000100110010101000110010100",
      "000101100100011001011000010000",
      "000010101001010101100101001010",
      "011111001101101001110101001110",
      "010101011000000110111111011101",
      "100001111101001010000101010111",
      "010111111101010011110010110100",
      "001101000100101000001100010010",
      "101011011011000100100100001001",
      "110111011011101001010111010000",
      "101111000010110111011100101011",
      "111100001110010010000101101001",
      "111001100001110100000001100100",
      "100100101101000011000100011111",
      "100001111111011000001010100011",
      "100000011001100001010010110101",
      "011100000011010110110000010100",
      "100000101000101001100101010000",
      "000100011111011111110011110000",
      "001101011011011110001100110001",
      "010000001010101111100101010010",
      "111010000010011110101111000101",
      "110101011110110101000101101011",
      "110000100011000111000101010001",
      "101010001010110101100000000010",
      "000101101100101111100111001101",
      "100110111100000011110000000001",
      "011110011100110110110011011001",
      "101000011000101101100110001100",
      "111011110101001100011100101100",
      "010000010101001100101011001111",
      "100110011100011110011000001001",
      "101100100100000111100011110011",
      "100100110110110110111100010100",
      "111010000010011001000011110010",
      "011001110010100000001100001011",
      "110110001011110011101000010100",
      "101110000110011100010101000101",
      "010001010000001111100011011011",
      "110010100111111110101001111000",
      "111001100100110000011000011110",
      "100010111001100001110110010011",
      "001010110101110011101101100001",
      "100110010001000110011010111100",
      "001010000010000110001100000111",
      "111011100111010100100000010000",
      "011100101100001011000111100010",
      "000011111101001111010101100011",
      "100110011001100101011011010101",
      "111000010110101110011110100100",
      "000110000100000101101110100111",
      "010011100101000001111101110110",
      "111011101111100110000011101011",
      "110110011010011100011010011101",
      "110011101100000000011100101111",
      "111000011111010010001100001011",
      "101010010000111010000101011000",
      "110001100111000011100110010100",
      "111110000101111110011101100101",
      "101000100101000000110000100110",
      "010011011011100111101100001001",
      "101101111111000011100001111101",
      "101000000010001101110011011100",
      "111001010100001010001101011010",
      "011001010000011001001001101110",
      "001100110100101000010101011100",
      "101011110000101011110101010111",
      "100010001010011010001000100010",
      "101000000100001100000001000000",
      "001111101000110011000011101111",
      "001110110011100011000111000110",
      "111000111101100000010001001010",
      "110001111000011011100000100110",
      "010110100100011111110010001000",
      "101000101100101011110111010110",
      "000100000101010011101001010110",
      "101101100000100000111010100101",
      "010100011101001011010010000101",
      "000000100011110011001110000100",
      "000100001111101110101111110101",
      "111001010000011110111110000100",
      "100011011110010110111001000011",
      "011010110110010011110001100011",
      "010100100110000111101011010001",
      "111000010000101101010111011001",
      "011100011101110001111001011000",
      "000010101001001011111101011000",
      "110111010001001101011011000011",
      "101001110110110101101110110101",
      "110101100110010101001111010001",
      "110010100000000111100110001011",
      "111001001010001111010100011101",
      "110110101010010110000011101000",
      "000001010011011110010111100011",
      "110100101001011010000110000011",
      "110010110100100101010011101011",
      "111011101010111111100000111001",
      "000000011000101011100001100011",
      "000100100100010111101001111110",
      "110000001001110111000100000010",
      "011001110011001100011101001100",
      "001010000011100110101100110000",
      "101011010000100100100010001011",
      "110000010100110101001100110000",
      "011001011010001110110011111111",
      "111110010001101101001100000111",
      "000110000100111001100100100001",
      "001010001001011100110000000100",
      "100111011010001000010010011100",
      "110110100000011001001001100011",
      "000001000011000000000010111100",
      "111011010101101110111111101000",
      "011000001100010000000111001101",
      "001010011100101101110100011000",
      "110000001010100111010001100100",
      "100011101111101000111101110011",
      "001000101110111001010011111101",
      "001010001001100111001011000010",
      "100111001110100000010111011100",
      "110101010111111011001111000000",
      "010111001010111110000111111101",
      "111000000110011100111011101101",
      "101000110110110011111100111100",
      "101111011101000000111001101111",
      "101011011100011100010000000010",
      "001001011010000001111010100101",
      "101110011111011100010001110001",
      "110111011100011001110111110111",
      "010100011010001011101100001100",
      "101111010011000001011111110010",
      "000011111110001101000111010111",
      "001111100001111111100111000101",
      "110101000001101000101011011111",
      "111011001001111110110101011100",
      "000011100100000110001001101101",
      "111111010001000011111010110011",
      "101110101001101011101001000110",
      "111101111110011011000001111100",
      "000001111000000110000010010011",
      "001111101000100000111011110000",
      "000010111100110011000011110110",
      "011011011100010011100110100001",
      "000110110100110110011010100011",
      "101110110110111101110101000001",
      "101001110110011010001111110010",
      "001100010011001110100110100110",
      "111001000010000110011101011111",
      "111101101101100001100010011010",
      "111000011001010000000011011010",
      "010001100110010110011110010110",
      "110001000111111011010000010011",
      "111111111011110011011100100011",
      "100000100110010101110111010001",
      "111011000000000000111010110010"
    ),
    (
      "001010100001011001010100111101",
      "011110111100101000110001000011",
      "010111011111110110110010011010",
      "011010100110101111001000010011",
      "110000011100101001011110001101",
      "001000100101111100010001000001",
      "100001110110011101000111000010",
      "010011100000011000111010001011",
      "110101001100001100111101100001",
      "100011101110101110011011000100",
      "010100100010100011110001000100",
      "110010010111110011010100001100",
      "011011111010000111110101110100",
      "101110110000000101110001101011",
      "111011100110111010001010000001",
      "110001110011111110100111000101",
      "110101000000101100100111000010",
      "010110000101101011100100010101",
      "100000110010011110100011011001",
      "111010001000011110111001010101",
      "110110100011111001010010110011",
      "000010011100011101010101001011",
      "101111000011000011010101101100",
      "001010011101110100111011110011",
      "001001010000011100001001010010",
      "110100111101011111111111110000",
      "011000100001110111010111100001",
      "010101101011000100001110000000",
      "011111011110000110100011011101",
      "110100000111101001000010100001",
      "010101101100001010011010001000",
      "110101001001110000010001010001",
      "100110101000010011111111011000",
      "011111111010110100000000110000",
      "010110000111101001000000100110",
      "001110000001000010010101101000",
      "111001011111100010100000010001",
      "011010101100011100011100000011",
      "011010000001001011111001010110",
      "100010011101101111110000010100",
      "111111000111101110011111001001",
      "010110011010010010011101111001",
      "110001010111111011001100111111",
      "101111000111100010000100010110",
      "000101100110110111101110010100",
      "101000101100101110100000100110",
      "111111110100111111111000010000",
      "101101100100010001010110111010",
      "000011110101000001011110000001",
      "001111011000010110001100111100",
      "000010000110000100001010010010",
      "111101100001010000011110000111",
      "100011000010110111001111100111",
      "110110110101110100101000110000",
      "010100011111111100100111100001",
      "111111001001100111010011010110",
      "010110010101010011110001011100",
      "001010000111001000101110110000",
      "111011101111101111000101000110",
      "101100101111000111101010110011",
      "111110101100100110101001111111",
      "011111110101100111011010001111",
      "101100101000100000001111001110",
      "110001011110010000101111001110",
      "101101010001101000100100111001",
      "000110100011111100101011110000",
      "010010100111011001111111011111",
      "111110100001010000100010001000",
      "001101011001100110011000011000",
      "001100010010100101111111001010",
      "000000000101111011110001010110",
      "100011011010101111011011110000",
      "100111100011110101100100011010",
      "111110001110001010101010011000",
      "111011000010110000011101001111",
      "010111110100000010001000001000",
      "111011001000011111001110111101",
      "001010100001101101101100101101",
      "111011011100111100000010111001",
      "100111101111101110011000011000",
      "001000000100011000110100110011",
      "111111001110001001101011100110",
      "101111000100111110100011001110",
      "000110100001010010100110100101",
      "101001110000011100010111110110",
      "110000110011111001011110010101",
      "001111101001100011101110011000",
      "000011110111100111110110111011",
      "010110100000100011111100101000",
      "001010010000001010000011000010",
      "111011110001100000011000011011",
      "001110100111100001001001001001",
      "011101000010010011000101101111",
      "010100001110111000111011001111",
      "101011010001111111000100111101",
      "111011110110000111100101101011",
      "110111011101101011010011000001",
      "001010001100010111110100111001",
      "101100011111101111101011011100",
      "110011110001011001011001111110",
      "010101000000100111111101010101",
      "101011101000101010000111110000",
      "000100110101000001010101011001",
      "111011101101011100001110010111",
      "110111010001110101011001001000",
      "111011000100100010101000101111",
      "001101111011101101101010010000",
      "111101010110111000111001100011",
      "010100001101011111111000001111",
      "110000010111001101011000110001",
      "000010101101111011010001101100",
      "001110110110000110110101110100",
      "110010100100110000101111011000",
      "011101110111100111111000110001",
      "101000010001010000111011101100",
      "110100011000100110101100001111",
      "011100010110111011001110001101",
      "101110101110011001100010111000",
      "010101000110001011011101101000",
      "110001111111101100010110111111",
      "010010000010011000001010101101",
      "000000111010000111110001010001",
      "101000111011111011110110011110",
      "100110111101011110001100001011",
      "101111110011000101010111001101",
      "010100100000111011110101100101",
      "110001110001011001001101001110",
      "011011111101100100100110000101",
      "001011111111011111011100111010",
      "111001000000011100110111110100",
      "011000011001110100100100010011",
      "101100011001010101001101100000",
      "010001101100010101001111101111",
      "111101110111010001000110111110",
      "100111111001111000000111010011",
      "001111110110100101110100110100",
      "100111010110110010011000110001",
      "011110010111000000000011111110",
      "010100101001111110100110110100",
      "100000100111111010011111010101",
      "100100100000110111100110000101",
      "010001000101101101010110110011",
      "011101101101011000101011001000",
      "010100111111010110101110001010",
      "101100010110000101111011100001",
      "111100101011011000100101100100",
      "110010101101100110001000101101",
      "011111000011101100001010001010",
      "111110101001011001010111110001",
      "000001111001001110110010100000",
      "100110111100000110011111011110",
      "000000101000011000001101011100",
      "011001010010100101011000000000",
      "011001110001001011110001100011",
      "110001010101101011110010110110",
      "111010001010111101001100000000",
      "010001000110101000101100000000",
      "011010010110001000000001101101",
      "111111011010010101100001010111",
      "011001001111110000010100110111",
      "000111100000010101000000010001",
      "100010111010001111001101111010",
      "001101111110100101010100011111",
      "111001001110001010111100110110",
      "100110010111001110101100001100",
      "100110110111001001011100010111",
      "000010011110000000111010001000",
      "110110011001001001001101001100",
      "111001101010111101110010111001",
      "101010101111010011000111101001",
      "111110100101011000101110110010",
      "101101100101101111000110011010",
      "111111001111111011110010111001",
      "110000110101111001011110110001",
      "101000111101110111000100100010",
      "010000000000000001010001010010",
      "010000100101001101111101110111",
      "001100001101101000000011110001",
      "001111101101111100010101110010",
      "111010110111001110001110100001",
      "011111010011000000111010111000",
      "011011010010100010011100100011",
      "000101000010111111001101001001",
      "011000000000000010000110011000",
      "010001011111100100010000110011",
      "110100001101111111100011000011",
      "001111110101001100101010011011",
      "110000111110011000000100000101",
      "001110011111111111111111010010",
      "011001111000101110000010101011",
      "110100000000100111011011110101",
      "111100101011011100001010000101",
      "111100100110101111101010001001",
      "101101101010111101001110100001",
      "111000011100111110001000000000",
      "111111111001011000101110010100",
      "111011111010101101010111100100",
      "100111010101110010110111000000",
      "110011111101011000011101111001",
      "111111010110011010000101000001",
      "110010000010111111101010000100",
      "010011110000000111000100110111",
      "111111001100111110000001011000",
      "101111110111001101011001011100",
      "000111111011010101001100101111",
      "110101011010010100001011101111",
      "101101111010010010101010001001",
      "100111101011000010111010000000",
      "101000001101100001000011110000",
      "001011100011000001111001011011",
      "111000000110011001001110011001",
      "100001100011011110011001011011",
      "010111000101110111111101000011",
      "111111000101010101011111000101",
      "101001101100110111100111111000",
      "111101101011100000000100011010",
      "111101011000010011100000101100",
      "000010111100101000101000101010",
      "011101001011010000100111010010",
      "010111001001100111111001000010",
      "001010110000100101010001111110",
      "101011111011000011111110111010",
      "101000010101110001110000111010",
      "001000111100111101110111111110",
      "100001001100100100101111001000",
      "110111101110000111011011101000"
    ),
    (
      "111110110011111001011001101110",
      "000001111110101111001010011101",
      "000011111000101010110100001101",
      "101001011001110100000101100000",
      "111110110110000110010000100100",
      "100011111001100101101000111000",
      "000011001111010001000101010010",
      "100011101011001001110110010111",
      "000010111111010110110111101111",
      "101010001011111011001001000010",
      "010110011001101000010001010001",
      "100100110011111011011001100101",
      "001110100101000111011110110010",
      "111010001010100101001110101001",
      "100110111000000011111011010100",
      "000000101111000100011011111000",
      "001101110100100111010000111010",
      "010100101101001101110100111100",
      "101010010111000101011011011001",
      "011110110110001110011010000110",
      "011111100001001010001010111100",
      "001100100010000000101110000001",
      "101000101001110010111001010000",
      "001110011100100110000111111010",
      "011000101111110110010010100100",
      "111101000111010111100101011010",
      "111000100000000010111010111011",
      "100010110110010001001101011010",
      "101110100001001011100110011000",
      "111100010111100011000010000001",
      "101010100011000011101100111001",
      "011100111000010110000011011111",
      "111101111010111111000010010101",
      "110001110101011111001010110110",
      "010010110111110011001111001011",
      "111001101110111101101010010011",
      "100001011100000110000010110001",
      "000001000010000000110101001100",
      "011110001010110010011100000101",
      "110101010001010001000000101110",
      "111100111011010100010100010000",
      "100111110000110111111101000101",
      "001000110101110100001101011011",
      "011001100100001101100100000111",
      "001100101101101011000000000100",
      "010110010111101000110100011010",
      "111011101111011101010010011001",
      "111011001000101100001101010110",
      "000110000110101000000010010001",
      "111000011000110011101000111011",
      "011110010101101101101111000011",
      "111011100011110010100111000110",
      "010010011111100001111001000101",
      "011101000100101111111011001001",
      "110111110001101001011101100101",
      "101001010111100000110001100101",
      "000100111100100111100110000010",
      "011111000100000011010111000110",
      "111001001100110101111101110010",
      "000001101000101000100100111000",
      "101010100001110011101101100100",
      "110101001000001101110010001010",
      "110011001001100100011010110111",
      "100101100010000111101100110011",
      "100001100101010001010101111111",
      "000001110010110101001111111110",
      "001010001111101101001011001110",
      "001010110111011100001111000101",
      "000001101010101001111010000000",
      "011111001110011000111011011111",
      "110110100101101101111100010100",
      "101000111010100000010100100000",
      "001111111010001110100111001101",
      "010110000011101011011001100000",
      "101001100100110011101000101011",
      "111101111010111110100011111001",
      "010100111111001011010010011011",
      "101011001001110111101100110100",
      "001000011011100010111110100000",
      "110000110010000100000111101010",
      "101101111001000100100100111001",
      "000111110011010011100101011011",
      "011110000000011101010110111110",
      "101000001000110100011111110010",
      "001001000001011110001011111111",
      "000000111100100101000000001101",
      "101000001101101110011010001100",
      "010001110001100000100011110111",
      "111100010011001011001011000001",
      "111001011111011010110011000001",
      "100110100110110101001110000011",
      "100101101100000001110000010010",
      "100110001000111101100010001000",
      "001100110011011101011000100011",
      "100011110001111110011010111111",
      "100111000010010010111101000000",
      "010001000010011010001011110100",
      "110000001001011101011101011011",
      "101000100110110011000100011010",
      "010101100010110000100100111001",
      "111110100001110111010110110010",
      "001001110101101000111000010010",
      "101010101001001100110001001111",
      "110011000111001111001101100100",
      "111111101100010100010011011001",
      "000000010110111000000010110101",
      "110000000011001000011101001010",
      "001101100001001101100000000011",
      "010000110100010011011011001111",
      "110110010101101010010111000111",
      "110011110011011000111000011000",
      "110100000110101100100000000001",
      "101110110000111010010000010010",
      "110000101101000010110011000111",
      "011011010110011011100011100111",
      "010111000001110111011101101101",
      "100000100011100000100010100001",
      "000010101111111111111100101101",
      "011111101000110101111001001111",
      "001100101011100001000001000010",
      "101000100111100011110111111001",
      "011100100110000101000010111011",
      "111001000000111110110001100100",
      "111100010011101001101001100011",
      "101100101001011010110111010000",
      "100101011101010110011100001010",
      "010100110010000111100001011001",
      "101111100110000100101010001101",
      "011101001101010010111001110110",
      "001101010110110011110111101010",
      "001100001010111101011111101010",
      "100101111100010110111010101110",
      "110011010111011110101011110100",
      "001101100000111110011001110101",
      "001110010111110111001110010110",
      "010011101011011101011110011100",
      "000100011101110111001101000111",
      "010111101010111011001000101010",
      "111111010011001001011011100001",
      "100100110101000000010011000000",
      "010001100100110011000000111101",
      "101011101101000101011001111011",
      "010011101011110100100000000100",
      "010001100101001110010100110011",
      "010110001001011100011011011011",
      "010011001001000000001001011010",
      "111101010010011111010010001000",
      "101000001011011101010101101010",
      "111100101001111101100010101110",
      "011111100011100101000001111100",
      "011100000100010110111110000110",
      "100111101110111100110001101001",
      "011001100010001101010011110110",
      "001110101000111100000101110100",
      "000010110001010100010110101001",
      "011011101000000101111011111011",
      "110001101001110111001000001110",
      "111100111111101100100111101010",
      "111110110111001011010010001010",
      "010010001100000110011110000111",
      "010100110001111010100110101101",
      "001001111001010000000011100110",
      "111000000000100110010100010101",
      "111000111110110110010000110111",
      "000011001100000111010111010011",
      "001010011001111000000110000110",
      "101111110001010101111100110011",
      "011100010111011111110011110011",
      "101001100011101010100010000110",
      "011001010010010111010101111010",
      "100011001110010101000100111111",
      "011111110100110111101010001110",
      "100000001010010001100011000101",
      "011110010011111000011001000110",
      "111001011011101000111000000110",
      "001111110010000100011011100011",
      "100111110111000001001101101110",
      "001111111011001010110110001010",
      "110100011001110000111101101100",
      "010001011011101111110011000110",
      "100100111010010101011001000100",
      "000100001100100110101001010111",
      "101011100110001110100000110011",
      "111101100010000000001000100001",
      "011110010001101011100101111111",
      "111111101110110001011101101101",
      "010010010011110111111010110001",
      "100010000100100001101000110110",
      "110100001111000010111010101000",
      "100110110011010010110001100000",
      "001010110001100000000100111011",
      "111110010110000110110000100101",
      "101110010000100101100110111000",
      "001011001111111001011001000110",
      "101110100100000000111100101110",
      "100001000111100011000011111101",
      "001101011000000110101000010111",
      "100100010000001100000010111101",
      "010100111011011110100000011001",
      "110000001010111011110101001010",
      "100000101100110101010101100001",
      "011111011001010110000111111011",
      "101101111110011111010001111110",
      "100100110111011010010010000111",
      "011110111110011100000001000111",
      "011100001010001010111101101010",
      "111010010000000110101101011111",
      "010111010010111000100001011001",
      "011011010001100000110010111100",
      "100011111010101010001101011111",
      "100111110100101110111110001100",
      "010000011101001101111100111110",
      "101001101101100011001011100000",
      "011100010100111010101001111000",
      "101111100011011101001011101101",
      "010010111100100011111011110111",
      "010101011101010100101011111010",
      "110011101000110101110000110001",
      "100000001111110101111011110010",
      "011010010100011101111101110111",
      "111111101111000000001011011010",
      "111101101001101001000010100011",
      "001001110110100110010000010110",
      "110010010110100000010110010011",
      "001010001001011111011100000000",
      "111101100001101000111010001010"
    ),
    (
      "110111011011000010111010011001",
      "011100100110000110111111100101",
      "000101000110001000000110001010",
      "001011101111011000011011011100",
      "010011001001011010111000101010",
      "000111100001110011001111011000",
      "001010010111011110111000111010",
      "100101100100010011110010001101",
      "111111010110010101010110001100",
      "110010100011010110111000100101",
      "110010101110000011011111000111",
      "100000000111111000101100010100",
      "110100011110100000011000001011",
      "110010101111010110000101001101",
      "001101010000111010100001011110",
      "000011101001001001100100000101",
      "011000100111011100010010010000",
      "100100110010011101101001111000",
      "000110001111111000000001110000",
      "001001100011101100001110100000",
      "111111100111010111101010111011",
      "100000011010000001001011010010",
      "101011010010101010001111010010",
      "100001011100100001101111010101",
      "110001011101101101111101000000",
      "111010010001011101111000011111",
      "000010011001010011111000010010",
      "011110111000100000111111000011",
      "000000110100010111100101110001",
      "110111011001001100110101101100",
      "101111001111001001110111100000",
      "101110000010001111011110111000",
      "011110000000011110111000010001",
      "111100010110101111011100010010",
      "001001000101111010011110011100",
      "010110100011011111100101000111",
      "010101110101001101001001111000",
      "101101100011100101110111001001",
      "010011001110011100111110101000",
      "010000001101100001000101000100",
      "001011101001011111011010111100",
      "111111100010000011000101101010",
      "101011111001110101101001000011",
      "110101001101110101110111000000",
      "000000110110111111001101100111",
      "000101110010111001101110000011",
      "101101100100111110110101000111",
      "000101010110010100100000110011",
      "111011111000010110111100101010",
      "111111010101010110011001011110",
      "111010011110000100110100010110",
      "010011110101111111110001111101",
      "111001100111000001100111000011",
      "001110001001001000001100111111",
      "100010110000000010001100100010",
      "110110001000010100101011111110",
      "111010001111011001111110000110",
      "100010000001010111010100000000",
      "111010111100001100101011000010",
      "110010001101111111111110000110",
      "111110100000111111110000011001",
      "010010111001001001000000100000",
      "110000000111110010110111101100",
      "011011110011010110100110101000",
      "111100110010101100011011011110",
      "011110001001100100001111101110",
      "000001110001001111001000100101",
      "001010010011001100110000111101",
      "011101011011011011010100110111",
      "001111001000100110101110100101",
      "010110111011101110101000011001",
      "101010100101101000011100010001",
      "111010100011110111101001101000",
      "110011001010100001101110001000",
      "000011101010011101001111100110",
      "011011101110011000011011111110",
      "100001000010111000000010100111",
      "010001101010000000111101001111",
      "001010010011101111010000100100",
      "011100111110000100101001010101",
      "001111111101001010100101110000",
      "101001000100010110001001111001",
      "011001100100110001100010011000",
      "101100110111111011100011110101",
      "110000011101001001001000110011",
      "100001110110000011010110111101",
      "111111001101000011110101001000",
      "111001100000110111011100000100",
      "000010111100011000111000111110",
      "101101010100101000111000000110",
      "001011001101011010101110101111",
      "101001101001111010011011110011",
      "111000011101010101000010000101",
      "110010011110000100101010100010",
      "110010100010100110110000000010",
      "010110000000000001011100000000",
      "110011010000100011001111110000",
      "011010011011001111010100010010",
      "011111010111001000101101110101",
      "111000111101110101000010100110",
      "011001100100001100000011111110",
      "010100100101110111001100000110",
      "111000100111010100100111011011",
      "000000010000110010110100110011",
      "111110101110111001011110010101",
      "101000110001011100001100100010",
      "011000011100000101011010011111",
      "010000010001001110010111111111",
      "000101010101010000011000010101",
      "100001011010110101110100001101",
      "100100101011100110000100111000",
      "000111100001111111111100101110",
      "111111001101011100111100110100",
      "001111101010101101100110110111",
      "010011001100000011100101001110",
      "000011010011110101011111000000",
      "000100010100011001111111101101",
      "101001100001011001011010000001",
      "110101011001000010101011010110",
      "001111101101101111010110010000",
      "000110111100110011000111101111",
      "000100000010101011110010010110",
      "001110011001110001100011011111",
      "111001110110101101110100111101",
      "100000010100110100111111000100",
      "010000011111111100110010010000",
      "101011100101100011110011101010",
      "100110010100100001101100001010",
      "101000100111001010111110111000",
      "101001001011011110101011011100",
      "110001000111110011110001011000",
      "010001110100000101011101011001",
      "100000110100100011000011101000",
      "100110100110101000010101100000",
      "000111000111010110111111101100",
      "101101110000011101001010010000",
      "001001100101111100111001000001",
      "011011110110010100110101010111",
      "010110111110000010000000110000",
      "111111000001010100011001110110",
      "011010101101001111011011100000",
      "100111000011011011001010111001",
      "101001111100110011100001011001",
      "101111001010011101111011110111",
      "000000000000110100010001011010",
      "111110110111000110001011110010",
      "001101110010001101110111101001",
      "001011011011111100110110101011",
      "001000010010100111010101000000",
      "001001000001100000111100101110",
      "110000101110000010011100001000",
      "101111111001000110001000111001",
      "111000010000001111010101010110",
      "001011100111000000111111111111",
      "011000011101110100010101011110",
      "111001100100011100010001110001",
      "101100110001000010001110100101",
      "100111010010110011111111100000",
      "110111010111101011011011110011",
      "100001111001110110010010011101",
      "011100001010111110010000011111",
      "000010111000000111010001111001",
      "000100001000100011011101101100",
      "111000010011101011010011010111",
      "110011010111110111000101011010",
      "100100001011100100011111011110",
      "111011101011101000111100010000",
      "001111000001101010010111111010",
      "111101111111001100000110010110",
      "001110000110001010101110100110",
      "111101101111111110100011100000",
      "000111110011111010001101001000",
      "101100110100111111001001101110",
      "000011111100110110001100110100",
      "000011110010101001110001011100",
      "011111010110111100101100000101",
      "101100101000011010101101010010",
      "010110110110111011100000001101",
      "110111110100010011010001111001",
      "100011110010100000001000001010",
      "010001101010111101111000001010",
      "011100110111000111011110001100",
      "010011101010000111000011001000",
      "100111010011101010100011010010",
      "110000011001001101111100011010",
      "101001110111110100010101100110",
      "110100100010110110101111000010",
      "100110010110110001111001100111",
      "100110010100010100110010100000",
      "011010011111110111011000010001",
      "000111111000111010101010000100",
      "011011000110010110100011011111",
      "111001100100011001001001111011",
      "000011000111001111010110011100",
      "111001001000000000011001011100",
      "101100000011110011001011000101",
      "110110111011010101110001011010",
      "110111110100000000100001111000",
      "000010000101001001011001100110",
      "110010010111011111100000011011",
      "100111011011100101100110010111",
      "101111001101101001101011010010",
      "101001101110110011100101011111",
      "111001111110101010000011000001",
      "010000111111111110111100001110",
      "100010000100001110000010001100",
      "100000000110011101001100000101",
      "001000001111001011010001010101",
      "001010000110010011100001010101",
      "011111110110110101101100001000",
      "100011001001100101100000001010",
      "101011000100110001000110000000",
      "100111110001111011111001100101",
      "010100010000000011101010011010",
      "110111010010001001100100001100",
      "111011100101101111111100101111",
      "101010001010101111011111011001",
      "111100100110001110010011010000",
      "001010001110010101010000001010",
      "001101001000010101110000000111",
      "110111001100011010100011111111",
      "000000001001111001011111110101",
      "010110001011000011111001101111",
      "011110001011011100101001011100",
      "101011011101011100100111101100",
      "100010000011010010101011000100"
    ),
    (
      "011011001101001011001101011110",
      "100010010000010001101111010001",
      "101101010010111011000101010010",
      "000001110011001110001101000011",
      "101001100101001000111110101010",
      "010010011111101111001100110011",
      "010110010101001110010111110010",
      "110001010000101000001101011110",
      "000110110010111011001101100101",
      "011011000001110101011010100100",
      "101011100101010011000011000100",
      "000011000100011010100110111010",
      "101100111101100100010001111111",
      "010000001111111011001101100000",
      "001000010101101100001010010010",
      "110101011011111111111011011011",
      "111000010011000011000100001111",
      "011111110000011001001010101101",
      "000011111101010100000111110110",
      "011101011101101001001100101111",
      "100000110100001010011010111110",
      "101001011001001000011001010000",
      "101001101011110101000010010101",
      "110100100001011100110010110100",
      "111110010011010000100110011011",
      "110000100001010011011010110101",
      "110111000001010101111001011011",
      "010101011110011111111011000001",
      "010100100100101010010000110111",
      "011001111000110010000100011101",
      "111111111101001100110110011000",
      "101100000101001111100101000001",
      "100011110010010101001101010000",
      "101110100101111100011100101101",
      "010000101000101110111111101001",
      "001111000010110110001101001101",
      "101101100000001001100000000101",
      "011010110110101011110010010001",
      "011010001111110010101010101001",
      "100001111001110001111110010010",
      "110010100101111111011000111101",
      "100011010101110100000101111011",
      "010111111010101110001110101101",
      "100110100100100001001100101011",
      "101011010000111010111101000000",
      "110010010100000111010101100001",
      "000000100101001001000110011100",
      "101101000100000111100101110001",
      "011010000100111101101101111001",
      "101111000001110000010011000000",
      "101000000010011110010011101011",
      "101010100100011111110011011011",
      "111001101101001010010100000000",
      "001111110001001010000011010011",
      "000110110110100111101001001011",
      "110101010111100111110100000011",
      "011000000000110101010011111111",
      "101111111110000100100010010111",
      "111000110111011001101110100001",
      "011010110001000001000001011111",
      "010000111000001110011100011010",
      "100110100110100010100010001010",
      "001000000000101110111111110010",
      "001100100001000111001000011111",
      "111001111010111010100111110011",
      "111001110101001001010011101010",
      "001000101100000111111010100110",
      "011110011111011000110101001111",
      "101010111000100110011000010000",
      "111001101000000010100110101100",
      "111100001101101000101001110011",
      "100101111010000101110110001100",
      "110100010011000101100001100110",
      "101011110101000110001000111001",
      "000000010100010001111001101000",
      "100111001010001011001111011110",
      "100101011100111011001110110100",
      "101111110000010101100000101100",
      "011010011010110011010111111010",
      "000010111110110001011111010001",
      "101111001110011100100100011111",
      "100111110010111001110111010110",
      "101110011101000101011100100110",
      "110011101011001100101111011111",
      "110011001001000111100001011111",
      "000100111001111100000110010111",
      "100101111100010001001000000010",
      "101111111010100110010101011100",
      "111110000101001011111011100101",
      "100011000010101111010100000101",
      "110000001111000111100100001000",
      "001010000000101010011010101001",
      "101100101000001110010001011110",
      "011011011110001001100000001010",
      "011001111000100010111010010100",
      "010001010100000111011100111001",
      "110001101000111101101001100111",
      "110101001110011010010010110100",
      "010001100100101000110001001000",
      "100000101011011000101111100010",
      "001100110110001011001000011110",
      "111111111100101100100001100100",
      "100100111000010110010110110110",
      "000000110100011101000101100101",
      "101111000010101000000001111010",
      "101011011111100000001111111010",
      "101110001011000110010101111110",
      "011110001011000101010000110010",
      "000101111000010101111100110011",
      "111010010110101100011001101000",
      "110001111001100000100111100110",
      "111010000111000101111010100001",
      "001001101100101011110111110001",
      "011101000101110000100100110011",
      "110110011001001001100111011011",
      "010000100110101100110111011000",
      "111000000011110001001011100010",
      "111001001011001011111111011100",
      "001110111011110111010000010000",
      "111110101010001011011100100101",
      "000011001000000100101101101000",
      "001010010001100001100101010001",
      "001010000000000011100010000010",
      "011010000000000010100001100100",
      "000100101111111010010010011010",
      "000010001100001100111100000100",
      "001101000001110000111010101111",
      "010001100101100000010001101011",
      "100000100110100100100110110101",
      "010110110101100111001000010100",
      "011011111011011100000010010111",
      "000000101101001111011110110110",
      "010101011001110110100101101010",
      "101011111000011001010111111011",
      "101001110101011011011000000011",
      "010001110111000011011100111001",
      "101111011001110000010000101001",
      "101110010001001100001110110001",
      "010101000111110010100001101111",
      "100001010111110101101001111111",
      "001110010110111011100101001100",
      "010011011011101110010010010111",
      "010010100100100110000001010101",
      "101010001011101110011100101110",
      "001010011110010111000000011101",
      "001001001000110111001111100100",
      "011000110101011110011101111111",
      "111011111011101101011110111111",
      "001001111101000111001010011111",
      "101110010101100101110110110111",
      "011010001100101011010110010010",
      "100100110000000101001010011100",
      "110010100111100100010111001000",
      "000000011111010110011001000000",
      "100100111101001110001001101000",
      "010111110011000001111001100101",
      "100110101100000000010011000101",
      "101111001100101101010101111110",
      "100011111100110011111001110011",
      "101110100011100000000011110100",
      "011111011001101101011110111000",
      "010110101010110100001101100011",
      "111011000110101010101011001111",
      "100011011011100000110010001100",
      "000100010011101101110101001011",
      "001011101000111011111101010011",
      "100101101010110110110001010011",
      "111001101000101010010111111111",
      "111111010111010111111010110110",
      "101000101001010110100010100111",
      "001111011110110100100110011111",
      "000110011011111011100101100010",
      "100111010100101001100011110100",
      "000100111010000111000011000111",
      "111111011010011110000011111111",
      "100010001010111100000001100010",
      "111111111101000101010110101000",
      "001110111101100100111010001111",
      "110001011001001001010011100101",
      "010010100010011001110110100110",
      "010011001110101100000110100100",
      "100001010010110100000100000100",
      "110100001011110100101111100010",
      "101110001111010101000111110001",
      "101110001010000010001100000001",
      "101001001101000110100001100000",
      "011111001110011010010110100001",
      "001111001001000110110010001011",
      "111101110100010011111100000001",
      "010001101011100110010001010001",
      "101010100010000110100110110011",
      "000001000010110011010000001000",
      "110010100000110000101100110111",
      "110010011000010101001011001110",
      "000011110010100100011001001111",
      "100100111000100011000010101110",
      "000101010010110111000011101110",
      "010011100111111111110111010110",
      "010111010011110011000110111011",
      "011001110100011010000010100101",
      "100011101011101001001001011111",
      "110110010101001000111110101000",
      "100101111111000100000001000111",
      "011001110000110111101001000110",
      "101011110011111110110001110010",
      "010100101001010011001001000111",
      "011101010000100010001010011101",
      "100101100010110001001101001101",
      "010111000110000000101010100101",
      "100011010000010110011100000001",
      "000001100000010100001001100101",
      "011110001100000100010000001010",
      "000101110101101000001101100011",
      "111101110000010111101110100010",
      "001111010010011011111101000100",
      "000110100101001010010101101010",
      "001111111000010100110101011111",
      "000001100111111110000011111010",
      "110100011110001110110111101001",
      "011101100110000100000100111011",
      "110111001001111001011011001100",
      "000100000100011010000011101001",
      "000110000101011010011110010111",
      "000010011000010011000110110100",
      "010110001001010100101001000001",
      "010111111000100001000100011000"
    ),
    (
      "010011110011011000101110001100",
      "011000101101111111100100100111",
      "010110010111111001010111000010",
      "000111001000100010001110011100",
      "001001010110001100110010100111",
      "010011101000101001110010110100",
      "001010100010111111001010111110",
      "001010000000011011110100101111",
      "101011100101000011111001000000",
      "110111110100111001011010000011",
      "100000001111111110011110001001",
      "000101001101011001101100011000",
      "111001000100110000010110000101",
      "111010010000111010011001010010",
      "111001001101101010100111011110",
      "101000101100111011010011011000",
      "000011100111010111100011001111",
      "100111000010100111111101111110",
      "111111010111010111011101111011",
      "011111101111001000000001011001",
      "111010011100011010011011000101",
      "100010110101001100110001111111",
      "001010100110010010110001010101",
      "101101000001010101011111111000",
      "101110001000111100000110000001",
      "101001100001001100101000100010",
      "111101110100010001010111110110",
      "001001101000000111110001010001",
      "011001111101010111011001110011",
      "100100011011100111011101011100",
      "010100010111010100110110111001",
      "100100100011111100101011011001",
      "000000000110111101001001111110",
      "110100111100101001000110100011",
      "101110011110110011111010011110",
      "110011101001010011000000010011",
      "010100010101001101010101001101",
      "101100101010011010011011011100",
      "001101101001100010101010001101",
      "111100101100101110110100111100",
      "100111000110010000000100110110",
      "101100000110101010000110011011",
      "110100101111100111010011000011",
      "010010101111100110000101111111",
      "000011000000010100001010011100",
      "001110010001101110111110001000",
      "100111101100011010110111100010",
      "010100001001010000110110110110",
      "001010010000000000111100100011",
      "011101111010010000011000000010",
      "010011100111111000111010111000",
      "100011000000010101010111001101",
      "010000111011011000000100011001",
      "101010000010110001110111100111",
      "000111110011000011111001010001",
      "011100110001101000111001010000",
      "110101111001001101001101111010",
      "100011100010001100111100111111",
      "001010001011101111001000011001",
      "001001111000101101001101110101",
      "100010001110010001001101101010",
      "101110011001001101011110001111",
      "100110101010011110001110001001",
      "011111100011000000000001000010",
      "100111111010011000101001001101",
      "010000000001011001011111110110",
      "000000010101110010100001000100",
      "001000000010111010010000010100",
      "010110101011011000011001001010",
      "100100011101100100101101100010",
      "011001001111100011110010001001",
      "001101101011101101110000010001",
      "000010000010011010000000111001",
      "011110000101111001010111100101",
      "101111100001010110001110111001",
      "110110100000010111011000000100",
      "000100011110010101001011001110",
      "001010101101000101101010000101",
      "101110101101001101000111101100",
      "100001010100100110100100000101",
      "100001011011111111010011101100",
      "110001101011011000111100010110",
      "001010001100101001110011010111",
      "111110101001011010101111000110",
      "001100100101101101110111001010",
      "001111110011011101011010110110",
      "011101111100111101101011111110",
      "000011001011011000000110110011",
      "010101000111111101111001011010",
      "000001011100011011010011001001",
      "100111100010110111001110011111",
      "010001110001011011000110011010",
      "001001001111110110010110100110",
      "010110110000010010001000111001",
      "001100111101111011101001011100",
      "110000001111000010011000010000",
      "110101111000010011010010011110",
      "010100111011011101110101010101",
      "111101000000111011110010011110",
      "000110101100000100111110011101",
      "010100101001101101001111010011",
      "010100011101100100111010101111",
      "110101001100010101100100111011",
      "100011011100010100110101111010",
      "101100000010010011011011000000",
      "100110011110100000111110011100",
      "110011010001000010010001110111",
      "011101101011101110000010010100",
      "010001001001101101101100000100",
      "100000001111110101000100001111",
      "010100000011000010111110001011",
      "101000101100111111110111001010",
      "010001000111111111010011010000",
      "111110101101101001100110000000",
      "010000111010101001101011011000",
      "011100010011001000111010000100",
      "111100010100110011000111010001",
      "110101000100011011100010101000",
      "100110000111100110111100010110",
      "110000010000111101001000011101",
      "110110101001001111011010000111",
      "000100100010101000011011110001",
      "010010001001111100001100111110",
      "101001100000001100100110101111",
      "111001101010101011111110000101",
      "111000110100101001100010110100",
      "001100011011101101010010011010",
      "110000000111011111101000010110",
      "111101101100100100010010010001",
      "010011111011101110011011100001",
      "000110010010010011101001000101",
      "111010101010110011000100011001",
      "010101001100010010001101011101",
      "110000101001110000111111100011",
      "001110110000110010110100100111",
      "001101010101110011100011000010",
      "110110101001100111101000111001",
      "111011111100111000100110101010",
      "110010001100001100011000110001",
      "001011000111111010001000011111",
      "101111101101110010011010101111",
      "001111010001010001111110000011",
      "111001011000101110010001100011",
      "111011100010000001010010010110",
      "011001001011011111000010111110",
      "010010111100100011001111011111",
      "111010000010010110101101110001",
      "011001111110101111000110001010",
      "001000100010010101010110001101",
      "011101000010111100000111110111",
      "011110001100011011011110011101",
      "110000001100101111101100010000",
      "110110110001010101000010000001",
      "011111000100011011101101110011",
      "000000101011011001000001111110",
      "110011111110101100110001001011",
      "000100111100000010101110111001",
      "100011101011000000111000010111",
      "100010100011101100001100111100",
      "110011000111100100110110010110",
      "101001010010101001111111011010",
      "001111111001001110100000110100",
      "100110100110011011000010110111",
      "010001110100001110110010011100",
      "111101101101011110101001011111",
      "010101111000110011000000101001",
      "111000101001110100100011110100",
      "100101101010010110100111010011",
      "010010110101010011110001100100",
      "010101010110100100001000011011",
      "111001000000101100111100111011",
      "011011010010001000101111010000",
      "001101010111001100100011100010",
      "011100000110111101001010011011",
      "110000011000101000001001001010",
      "011101100100000000011011100100",
      "001100110101001001011111101100",
      "100000000111011001100111001110",
      "101010111110110011001111000111",
      "010110101100011010111101100000",
      "011100110100010001010001011001",
      "111011101010001101000011001100",
      "000011000101101000100001101001",
      "000001011011010010101001000000",
      "010000011001000011101011100000",
      "000001000111001001000000111110",
      "011111000100110111001001000011",
      "011011000100100010000110110110",
      "110001111001010100010001011001",
      "010010101110100101110100101001",
      "011000001110100011001110011100",
      "011000101011100101101011110110",
      "100010000000101101001001000001",
      "101000111110100001000100010000",
      "011110000000101011110011100110",
      "001000011011010101100011111111",
      "010010110000000000001010000110",
      "111100111011011111000011001000",
      "101011101110011000010011100011",
      "110111000001010000011101111000",
      "001101100001110000111001101000",
      "101111010110001011000110101010",
      "001010111010100001010011011100",
      "010110100000100000001101111111",
      "010000000110110101001000110010",
      "101001011000010100010001011001",
      "100111101000101100001011000100",
      "000000110010010100010101000010",
      "001010100111110111000100111110",
      "000111001111110111010001101011",
      "000101111011101111011010110011",
      "101101101011100011111011111001",
      "101111111110101101100100001000",
      "101000100100101001001011010111",
      "100110000110001011000101001010",
      "000111111010000000110101100010",
      "001101111011000011011000010101",
      "011000100111010110000100010101",
      "101101000010100000010111000110",
      "100010100110101010001001111101",
      "111111100000100001010001010001",
      "011100100110000111000000110101",
      "110011101100000100110111101010",
      "111010111110111001101011110001",
      "101001111010110110000110010100",
      "001000111001011011111011011010"
    ),
    (
      "001100010111100010011001110101",
      "011001001100111110110101111110",
      "101010101010100001010010001000",
      "011111111001000101011011100110",
      "110110000110111111101100110111",
      "000111011010010011111010110110",
      "101010001101111100110000011000",
      "001011001000111011011011000000",
      "110101000110111001001011000000",
      "111001110010000111110111010000",
      "001000101111000011011010010001",
      "011111111010100000101000000100",
      "001111110100000010000001111110",
      "110001111111100001010110110101",
      "100010101000010000010001001110",
      "110011110010001101010010011000",
      "100100000100101000100100011110",
      "011110010010000011110010000010",
      "001100010010001111001010111010",
      "001000110000010111101001000011",
      "011100101001111111110101010101",
      "010001100110110000000011010001",
      "011010000110111000111000111010",
      "011101011101111001100101000010",
      "001100001010100010000010111010",
      "010000100101100000011010011000",
      "111110011001101000010000110100",
      "110100101000110011111110011000",
      "100111110100001100000110100111",
      "000011111010101000001111000101",
      "000010001000101010111101001000",
      "100101011111010101100011010010",
      "101010001000100111100011001101",
      "101100001001010001010011010111",
      "110111110001111110101111100011",
      "010000101011100101110000010110",
      "101000001100110000010111101100",
      "000010011011001000100000000010",
      "000111101111010001110101101010",
      "000001011010111011110100100011",
      "111101100101011011111000100010",
      "011001010100010110001000100110",
      "111001010111011111000111001101",
      "001010110110100100011010011001",
      "101011011111101100000000000111",
      "110001111111000111001111111100",
      "110010010100010001100110111011",
      "110011011001010111001001000100",
      "000101110010001111001101100100",
      "111010010110011001011011100010",
      "010100010110111001110100110000",
      "001101011101011101110001011111",
      "000011011000100000101101011011",
      "001110010101000001000010110111",
      "011001001010101110000010011000",
      "101110000001011100010000100001",
      "101011001001111010010000000100",
      "011110001000010100000011011111",
      "001110100000111111100011000011",
      "010111100010010100101011111000",
      "101100010111010100010010011110",
      "101010011011100110001000000101",
      "010011100001010000000101110101",
      "010010101100101110100110010110",
      "001110111010110010111011011100",
      "001000100100011011010000000010",
      "010011111100100010111100100100",
      "100101110100111110101000001011",
      "001001001000010111110101110011",
      "000010111100001010110010000010",
      "111111100111011000110001101110",
      "001100100101011001100000010011",
      "000000111101001100010011101001",
      "010110011100111100101110000001",
      "000100011010000010100010111100",
      "011100001111110100100011101011",
      "011111111010110101110110110111",
      "101111100000000010010011101100",
      "011101010011000101001100101011",
      "010111010010110010011010010011",
      "011000111100010111000111011000",
      "010100110011011100000000011110",
      "011101100010100100101100101010",
      "011001001101001001111111011000",
      "100111101101011011110000101001",
      "011001110100101010001101100011",
      "010001011111110010111010011110",
      "101011011100010110011001000000",
      "110000000111011010111110011010",
      "110000101111010101010010111101",
      "111000011100101110110011111011",
      "001100000100100001100001011011",
      "000001111000001010101000010001",
      "100001011101011001011001101010",
      "110011001111011110111011001110",
      "000110000011111101001111101110",
      "001110111010100111000110100111",
      "000110111110001011101011101001",
      "110100100011011101011011100001",
      "101001010101010001000110001001",
      "010011111101011010111010110001",
      "011111110111010110101111110110",
      "100101001011010110101100001000",
      "001010011010000010000011110001",
      "110000101100100111110011001010",
      "010010110101010001000100010010",
      "100100011101001101010011011000",
      "000010010010000000110000001001",
      "000100111111011100000111111110",
      "101111101100001011001010000000",
      "000001110111001010101101100010",
      "011100000110100110000010111001",
      "100110001111000011000110100110",
      "010111010000011111110010110001",
      "100011100101000000001000100001",
      "001101001101100100110111011001",
      "101111111010010101001011011011",
      "000011010101100000111001000110",
      "100001100010100011101001010110",
      "111000011110101101100011011100",
      "111101101110110011100011110010",
      "110111111011101111001111001001",
      "011100111011001000000100111001",
      "000100100111101111110111100011",
      "110100100110001010101110010001",
      "011000001010110100100000000111",
      "000110011110000101011001111111",
      "001001011011101001100100110100",
      "011101000011101011110011111000",
      "010110011011011010101110010000",
      "010111011001100100000100010111",
      "000001010110010000111100010010",
      "100111111100101010100011010101",
      "011001011001010110100101111001",
      "110000001111000111000001010111",
      "101100101110101001111101001000",
      "111100110010101001100011101100",
      "100100000111010110011101101111",
      "100001011101001000000011101010",
      "101010010001001101001110000110",
      "011000100100000010010101001000",
      "001110000100100001001110000011",
      "100110011101010011000010010111",
      "100000010111000110011001011000",
      "011010111100100111100010110000",
      "111111000110010010000111111111",
      "111110100101111111010001111100",
      "111000011100110011101100000100",
      "100111011101001110010111111011",
      "011000101100110110001110001001",
      "001110011001110101101111110000",
      "110100011000110010000011010011",
      "011011100010110000011111011001",
      "010001010001001011000100110110",
      "010100111001001110011110001101",
      "110000101100000110110010011001",
      "100011000100111100100100010100",
      "010110010110110000000010011100",
      "100100010011000111010010011001",
      "101000001000111000111000011110",
      "101000111110101101000100000011",
      "001100001100100011111101111100",
      "010100111011101001101010111101",
      "000110110000110101010010000011",
      "110000010101011100011000100001",
      "111110111000011001000011111001",
      "100001111111110100101101011110",
      "011001101011001011011011000001",
      "010011001100110110111010001110",
      "000010001000111100101111011000",
      "000011110100010110101010100110",
      "101100110001101100110101101011",
      "000100000001001010011101111000",
      "000011110110110000110111001000",
      "111110111111110100110010110011",
      "001100111000100000100011010101",
      "110000101110010111001101110011",
      "011101011010111110010101000101",
      "000010000101001100001111000000",
      "001000001100010111111010101101",
      "010110011101010001100101000011",
      "011101110011101100011100010001",
      "111101011001000101001111101100",
      "110000011000000101000101101100",
      "010100111111111010001001011100",
      "100000011110100010111010001001",
      "010111000100010111110101101100",
      "111000000001110110010010000100",
      "010110000111001001010011000001",
      "110111011001000001110110110101",
      "100001101001111111100100100010",
      "111111000000111001110000010110",
      "000000100111101110111111110011",
      "101111011011110110000110011100",
      "110100000110100010111001100000",
      "100101011110000010011010010111",
      "100010100111101000001100111001",
      "110010010011110101010010110100",
      "100000000001001000000011010110",
      "101010001101001110011100111110",
      "011001111000010100001000100101",
      "010111111001011101110010111100",
      "001011100100101111011011010010",
      "000100100001000101111001010010",
      "011100101110111100000011111100",
      "100111110111110101011100000101",
      "000000100111001000101100111101",
      "011100110011011110000011101000",
      "100010011101000100001000000001",
      "010100101100110000011011011111",
      "011111001001110011010011000011",
      "010101001101110010101110010111",
      "000101010001011110111100010101",
      "100111011111101001010010111011",
      "001100000011100101100100000001",
      "010000111010001100111101111010",
      "001101110010111001010010011101",
      "000001000110101010000100110010",
      "001010011100110110101100011101",
      "011110110100011011001101010110",
      "011011110110110110011111110110",
      "011010100011000001011100100101",
      "111001100001110010101110011000",
      "110000010111101010110000000111",
      "000101100000100110001011110100",
      "111011111001110100110001001111"
    ),
    (
      "010011010100010111010101111010",
      "010110000010110011000111111001",
      "110110011100110011001110011010",
      "011111000111011000011001111100",
      "001110000010010011001101100110",
      "001010110010110110000101001111",
      "000100100010001111101010100100",
      "001111000111000100100100001100",
      "001101111010101010101100011011",
      "100110010100010111101011100001",
      "011000011111010010010110000001",
      "101100111000001011011100000110",
      "011101000101110011110100100101",
      "110110110001000010101100111001",
      "111111110010000000100000101010",
      "000100110011110000101111010101",
      "110011000010001111000011000101",
      "100101100111001000010100100001",
      "000010011101101111010001000001",
      "001010010011110001000011111001",
      "100101011110101011101001011011",
      "011001001000000011100010001111",
      "101111000110010010100010001111",
      "101100100011100100111001111001",
      "001111110100011111110110111111",
      "111110000001111111101001100111",
      "000010110111111001110000101001",
      "110111111110101000101001000010",
      "110100010111100101100110111101",
      "011001011001101001110111111000",
      "010100100110100010001010111010",
      "111110011110111111011100111011",
      "010111001110010101001001000011",
      "010100100101010011111000001101",
      "010101110110100101010110010101",
      "001100001111000001100101011111",
      "001101101100011001000110100111",
      "100101101010101110011110101101",
      "010111001100001000000000111110",
      "100010000100101100011001001000",
      "110000000111111111111110100101",
      "110110110110101101100101110010",
      "110011000001111111001001111110",
      "101100001001100110100111111010",
      "011000110101000101110001111010",
      "111001010111101101000111110000",
      "101011001000110101011100000011",
      "010110000100110001001101011001",
      "111011000110111000001100101011",
      "110100001101010000001010011011",
      "111001110000111110111110111000",
      "100000101011101101010000111011",
      "111110111111111110100000010011",
      "111101001101101100111001000101",
      "000000001010111111101111101011",
      "010101111100110010001101011011",
      "010011110101110100110100010011",
      "000110110100011010111100100001",
      "111111000001001001100101011100",
      "011101111100110110000110101001",
      "110010101010101000011000011111",
      "110001110000101110010110100110",
      "110000101001111110010010001010",
      "111110000001111110111000001100",
      "100100010000101011011001001011",
      "011101010111000000101011011010",
      "011101110000100011001001110100",
      "111110101110011011110000111010",
      "110101111010100011111100001110",
      "001001011011011011100111110001",
      "000111111111011100000000010110",
      "101010010001010010010000110100",
      "011001010111110101101010110010",
      "110101101000000110100101011011",
      "100011001001010100111010110000",
      "110111110101100010110010010000",
      "010100100010001001011011100001",
      "101001010101011001100011101100",
      "001111100000011000010111100010",
      "001111010011010110010011110100",
      "100111110011101100000100010110",
      "000010111001001101110001111111",
      "010001001100101110000111111011",
      "010101110100110001111010110001",
      "101111111100111001000111011100",
      "001100000001000000000001000100",
      "100011111111111101111110110100",
      "011101010110100100111111111110",
      "100100110000100100011011011101",
      "101110101110100101000111100000",
      "001001010010111000111010111000",
      "000011111001111101110110110100",
      "001000001010010111011010001110",
      "001110001101000101110111110011",
      "100001100111010100110011100100",
      "000000000111100110101101111011",
      "010110011010010111001000100110",
      "110110100011100111001001101001",
      "010111001111001001100100100100",
      "101100100011111111011101101110",
      "010111101011011001111010100101",
      "100001110100011011011101001100",
      "001000110111110000010101101110",
      "011101101100110101010000010001",
      "110100010011101001101010110110",
      "011010011001111001100111100110",
      "100000001101111111111101000011",
      "010110101011010000001111101100",
      "011100101101101111000000000010",
      "010010101100110001101110010100",
      "001100001110101000000110011000",
      "100111001101111000011000101101",
      "100111001100101011000010011100",
      "100010000010101010110011001111",
      "101011101010101111010110100001",
      "111010011011011111100001110000",
      "000111001110110100110010000001",
      "111111111010011101100010111110",
      "000011010101010110001100011100",
      "100100101110011000001011111011",
      "100000001110111111011110010001",
      "011010110100100110100001000010",
      "101111100010110100101000010111",
      "000100000101100111001100110011",
      "100110101010011010111110001101",
      "111011101011111111010110010110",
      "101100011100001101111100000011",
      "010001110111010011001001110001",
      "110110011000000010001101010111",
      "010000011101111100100011111100",
      "111011101111010010010011010001",
      "000100011000101101000100010000",
      "111011000000100111000111101011",
      "101010000111110010010000101100",
      "000000001011111100101110001010",
      "110110010101101100011111010110",
      "001111100000010100010111101000",
      "000011010010010110011101011110",
      "001010100000001111001100000101",
      "110110010111010000010001100011",
      "011111110111011101000010011001",
      "000100001101000100100011010110",
      "110001011110001100100011100000",
      "001111010100001101000111101010",
      "110001110000101010110101010100",
      "110010011010100111100111111001",
      "111011101100110011110101110010",
      "101000100111011100010101011100",
      "110111111111000101010000011111",
      "001000101011110100111000001000",
      "000011100100010010011100111000",
      "101000101011111010001000111011",
      "001110101110011111101001001000",
      "001000100011010110110010101000",
      "111001101011000111111001111011",
      "000111101010000100001101001110",
      "101100100011001100111111011000",
      "010101101010000010101111101100",
      "001000100010111000011100101101",
      "010100001000010011001011101000",
      "110001011111111011011101000100",
      "000101100001100101101100010000",
      "001000101011101011000000100011",
      "110101111100001010000111010101",
      "110010010110110010010111010100",
      "110100100001100101100110010111",
      "100100000010101101010000001101",
      "111000011101011101111100010101",
      "110111010010110000010001010011",
      "011011110110101011110000101111",
      "110100011101010110110110101101",
      "011110001101010000110111110001",
      "111101001101101011011010100100",
      "011011001110000011111111011110",
      "001011001000111100011100110110",
      "000100000111000111010000110001",
      "010010000110111111100000000011",
      "111000110001000111000000110001",
      "011000110010000100110001100101",
      "111001100101010100110110000010",
      "111110011111100110111010001011",
      "111001101101011010110001101001",
      "111011001001111011001011010111",
      "001101101010101100110100100111",
      "110110110100010011110101111101",
      "000011101100011100010100010110",
      "011011001011001101001000111000",
      "010100000110010000010111010011",
      "001101010011111000101001111001",
      "101011010101011110001100001101",
      "110010011101101001000011000100",
      "010100100000100010100100000001",
      "100011011011001111011010110110",
      "101111010011010100011000000110",
      "000111011111110110010101101000",
      "101101110001100111100001001000",
      "101111010010010101010110010101",
      "110000101001101001011010110011",
      "101010101000001000100101110001",
      "100010000001000011111111110100",
      "000111100110010010100011011110",
      "111101010001110100010100111100",
      "000101101000101001001100110001",
      "100001010001101100111110010000",
      "000110001010110001010111110011",
      "100010101110010110111110111001",
      "011111000110011011101110110111",
      "101100010000100101111101010000",
      "001001100110000101011110110100",
      "011110100111011110000110000111",
      "011000110011010000101111011001",
      "100100101110000111001111111110",
      "011110011101101011000110101111",
      "101001011000101101010111100100",
      "010101001000001110011110010011",
      "001000011110010000011100000110",
      "010010111101111001010101001000",
      "100110100001111011011101111001",
      "000111101011010101111000000011",
      "011111010101111100000101111100",
      "010110110001000100010011011000",
      "110001100000010111111110100111",
      "011001110110110010001010011101",
      "010010001110001110000001111010",
      "110110011011111000010110010000",
      "001010001011011110001101000000"
    ),
    (
      "101000010110101110011011011110",
      "000100001100010111001101110110",
      "110010010011001010100110110000",
      "101000111111011101110011011011",
      "100111101000011101111010110010",
      "000101111011101100001000110101",
      "110101101010000111001001001111",
      "100011111001100000000001001010",
      "010010111000011001001111110010",
      "100101110110100100100100010011",
      "011001001100010101011110101101",
      "101101100011101111110101111011",
      "110100011110100111110110001010",
      "011110000001111100101101101011",
      "111011000001111000110011111110",
      "111100111100010100100111000000",
      "001100101101111101010000110001",
      "010001011110101101010010001011",
      "111111011101111011111110100011",
      "000010011111110010011110101110",
      "111011000000011010011111010001",
      "000101101000010111011111010011",
      "111100110000101101100100110010",
      "101101011110011000001011010110",
      "110101010010110111111101110001",
      "001111101111010101101100100111",
      "000111010100000100000000111111",
      "011000101001101001101100001100",
      "101011111011001110100111111011",
      "110101111001101100001100010110",
      "001001111011110011000011000110",
      "011101011011011101010101000011",
      "111101000001011010001001111001",
      "011000010001101001111100101101",
      "011001001000001110001110101000",
      "110011110011110001001101010101",
      "001110011100111010010110110101",
      "100011110101101011101001100110",
      "110000010001001011000110011000",
      "011110111000100010011110100010",
      "000010110011011010100011101011",
      "111001110110000111101101010110",
      "010011010111000101110100001011",
      "010001001011110111001101100001",
      "010110101111000001100110001000",
      "011010011100001000110100101101",
      "000101110011101100100111100000",
      "110101010100000101010101010011",
      "001101001100100110001001101011",
      "010100010111111010000111110111",
      "111101110101110011101111001101",
      "011001101001110010101001011110",
      "010001001010011011010010101011",
      "000110101101110011100011101101",
      "110100000100001100101011101010",
      "101100000010111010010010110100",
      "001000100111000010101101010010",
      "001000100001111000000011111100",
      "111100010010000100000101001011",
      "101010101101110111101101111000",
      "100001101010011000011111000111",
      "011010100001010001000001010110",
      "000101001101011011111001101110",
      "110101111000001110101101010100",
      "110001011011101001111001110111",
      "011010010010101001001101100010",
      "000011001011110011100000001010",
      "011110010010011100011110001000",
      "101010011011000010011110110011",
      "011110001101101101101000001100",
      "010101001000011111000000000111",
      "001011000010010111100010101110",
      "011110010010111000001001111010",
      "111000110010111111101001101110",
      "011001110000000011111100110001",
      "100100101001000101100001000110",
      "110111011101011001101010110000",
      "000011111000001010111101000011",
      "110110111101101011001010001010",
      "001011010010100101001000000101",
      "010001010001001011000000101010",
      "101110000110111001111110000111",
      "011011000110010100111101000100",
      "101100100010011110100100100010",
      "101010110001010010000101111111",
      "110010011010000011001011100111",
      "001010111110100101001000010110",
      "010100000110110111110010101111",
      "000101000111101111110000000000",
      "010011001001111010000010111101",
      "100011110111011111101110110010",
      "101001011100111110001101111101",
      "010111100101101011001000101000",
      "101111010101001100011111111101",
      "111100000101011101000001000101",
      "001011110011010100001000101001",
      "011101110001010011101100111010",
      "001101010011011110000000101011",
      "011010101110111000100110100010",
      "010101000101110010000110001010",
      "111110000011111101001100000010",
      "111111011111010001011111010100",
      "101001001000000110100000101101",
      "000101010100011000101110101100",
      "111011000011001010101101111001",
      "100010100010111111110011111000",
      "010100000101110101001001111011",
      "111100001011101010001000011000",
      "010001100111000111111101111110",
      "010000010010010111000000111101",
      "110101001100111110100001001101",
      "001101000111100100001101011010",
      "101101011001010011110010100101",
      "101101101011111000000001001101",
      "111100101110111100001000010001",
      "111111110110111111110101101000",
      "111001110011101001100100010110",
      "000010111000101111100110001010",
      "000100011100001001110010110100",
      "000100111100010000110111001000",
      "001110011010010000101110111110",
      "011110111011111010101110110011",
      "100110001101000111000110000011",
      "101000100000110111000010001011",
      "011000011100001000111110011100",
      "110101110101001110100011101110",
      "101011010000101111011011101110",
      "010111100011101000000100101010",
      "111101001110100110000001000011",
      "111010001100011011010111101010",
      "100111100101100100001011011111",
      "011010000000101010101111101111",
      "101011111011000010010111111001",
      "101110110101011101000101111000",
      "011100011001100111001001001001",
      "011111001000000001110100110010",
      "011101011110000101011001011001",
      "001010000111101111101011001101",
      "001001101101101101100101010100",
      "011101011100011111011110001000",
      "111011010101111110001010001001",
      "101100110010100100000111101010",
      "100100110110001001111010000000",
      "001100101101111101000000000010",
      "010110000000001011101010101101",
      "001010010101101110000111110010",
      "110001110100001010001101010001",
      "010100000101000101010000100001",
      "101111000111010000010000000101",
      "001000011001110100000000110010",
      "100010100100010000111110100100",
      "101000101010001011100101010110",
      "101111010110111001100001110110",
      "101111101000011111000000101011",
      "100001011011000011000101000010",
      "001001000110011100011111110000",
      "100100011000010111011100001011",
      "001010110100000111111000111011",
      "100011110100011110100000000110",
      "110000101010000101100111101101",
      "000011101011010111110110011100",
      "001110110111101101011010110011",
      "111110111000001000000000001101",
      "011101011100101011110111111010",
      "011101110110111110011011101000",
      "000110100000111000001010101110",
      "100000101110001001011100100000",
      "110011100101110100100110111100",
      "011111011010100001010010011100",
      "100101111010101001011110001101",
      "100100011000110110110100111110",
      "011000101110111001011110101010",
      "000001011010010111101001101011",
      "011100101110010010000100110111",
      "111101100101101001000001100001",
      "010110011011101011010111001100",
      "010010010000011110010011000100",
      "001001100110001010010111101010",
      "100011100011110110111100000111",
      "000000100000000111101000010001",
      "110010101000001110011101110100",
      "110111101000000010011010101110",
      "010110000111110000001110011110",
      "001110011100010000101111001000",
      "000001100011101001001101000010",
      "101111100000101001110001100110",
      "110010011010001101110000101011",
      "111101100000100100101101110100",
      "010011001100001000110110011000",
      "001101111011111110000110100110",
      "000011001000100111110111100100",
      "111111000011010100100111011000",
      "111111100000000111111011000000",
      "111001001101001000000100010001",
      "000110101100100010111111000100",
      "110111110000111100011000011110",
      "011010111011000011010011100001",
      "111010100001010001111110110000",
      "011111101001100111001000101000",
      "000000000000111110101000011101",
      "111110000101100110000011101110",
      "110000011001110101111110001101",
      "100011010001110101101111000111",
      "101101110001110011001010100000",
      "100100000011110111010010010101",
      "101100110101011000100111011101",
      "011101011001110010011011001000",
      "011000101110111010101110110100",
      "011010101000010111010111111111",
      "010000010001110000000100100000",
      "101110010011101101101101111011",
      "010111101100001101010110001110",
      "100011111010110001011101001011",
      "110000001000011010011111111001",
      "101101001110111000101110000100",
      "000010010010100101100011111100",
      "001101011110101001001100010000",
      "100010111101100111001110111110",
      "010110010001101100110001110011",
      "100010011001111011011110000001",
      "001000101111111000000001100101",
      "010001011001000011000011000111",
      "100100001111101110001000101011",
      "100110001110101001100101010110",
      "000000000110000101001110111110",
      "100101100010010100101101110100"
    ),
    (
      "001101100110000101011101010111",
      "100110010111010100000001001000",
      "101110000010101110110111101110",
      "100001100010111101110011011111",
      "110101010001110110010100110110",
      "010001000100101000001101011111",
      "111101100000101111000100000010",
      "000110000110010011110000010010",
      "001101010001100110001011010100",
      "111100101011010101111111000110",
      "101011101001111011100100000010",
      "010100000011110111011110100001",
      "011111010101110110011011010101",
      "001100101010001101100010110100",
      "100110001110000000100000111111",
      "011010011010110000111010010000",
      "010000000110100000101011110100",
      "001011010110101001101010000100",
      "001000110110110010001111100100",
      "001010111001001101100100101111",
      "110111001000000100010011101011",
      "101101010110010001110100000001",
      "011110111111000110111010101011",
      "010000010000011101000111010111",
      "101111101111111001000010111010",
      "010000100110001000000011111111",
      "001011010100101101101111000110",
      "111000011000111001110100001000",
      "110010100001110011110000111001",
      "011101101010101010111000111101",
      "101000010010100010011001100001",
      "001100110000010110010010000110",
      "011111110111101111011001100011",
      "001010101100010111011001010000",
      "110100001101100001000001100100",
      "101011111011010111001001011101",
      "110001000000011110000100110101",
      "011100110100100010011000111110",
      "101001000101001111111001000110",
      "110110111000001001010110010000",
      "110011000010011101111101111111",
      "010011001000100011110101010011",
      "101011010111111001100010000110",
      "010110110110110010010001111110",
      "010010001011011000110110110011",
      "100111111001100110010101100001",
      "000011000110011110000101001001",
      "001100010100000100010111100010",
      "001001110011101100101000110110",
      "011001101010100100000000011110",
      "111111011101010111100010101100",
      "011011101110010100100110010001",
      "111110001010000110110111100001",
      "011110001000011111110010001110",
      "100010011100101000110011000111",
      "111101001000101110001011111101",
      "101010100000010011000000000001",
      "101011000010101011100001001011",
      "001110110101111001101000101011",
      "001101010001010000001010111011",
      "000111010101111101011110010101",
      "101110001010111110001100111001",
      "001011011110010010100111110101",
      "100010010101111110011000000111",
      "010010000101111110111110000110",
      "001000111101100110011101001000",
      "010001001001010100010011111101",
      "000011001010101111111101011100",
      "111111101010100001110110001001",
      "011001111110101100101000101001",
      "010100001010110001101101011110",
      "010101110100010011001110110010",
      "111011110001111010011101001000",
      "111000010111011100010111010110",
      "110111001101001001001010111111",
      "111111011000100010111000001010",
      "101011010111111111001100111001",
      "001011110010100010000110011110",
      "111000110101111101101110010101",
      "010111110000101000101101001111",
      "101011010001010011001010000101",
      "001000100100000010011000001111",
      "100101001000010011000111111001",
      "011001110111000010100010010101",
      "010101010100011001011001010111",
      "001110010001100111011010110001",
      "010110001011000001001110000100",
      "100110011011011000000110011010",
      "110001001101000100000001100100",
      "010110100111101101010100011010",
      "010110111001011111010110110111",
      "001001000100000000111100010100",
      "010001111000001001000101001000",
      "100010110010110010111111100000",
      "011000111011001001100010010000",
      "000110001001011010100000110011",
      "110011110101111011011110101001",
      "110111001001100100110001101010",
      "111110011110011100110101100001",
      "011110101001101111001000101100",
      "100100000100011100011001110100",
      "000100000010100110011100101000",
      "111101010001010110111111111110",
      "101100111010011000000010010100",
      "001110010010001001011111011110",
      "010001010011011101111110001111",
      "001100000000100100001100011010",
      "011100111010001010011001111100",
      "011000100110100011101011010001",
      "000110000010011001010000010010",
      "101101110000101001010010001101",
      "111000001111111011100111000100",
      "000100110000110111100111110001",
      "111010100011100100001100010110",
      "101000100100111111100110101011",
      "100011100001100111001011000010",
      "110101010110101110010011011101",
      "100011110011100101100111011110",
      "100001001101011111011111010011",
      "001100001000011011011010111101",
      "001010100000010110110001111011",
      "101110011001111010001001100011",
      "000110010011101011100000110000",
      "100111010010000101011111101110",
      "110011111001110001001100111101",
      "000110101101011011100010011100",
      "011101000010011110010001000000",
      "010011001111010100110011000010",
      "011010001010111011000001001011",
      "111000111011011001101011111100",
      "101100001110010000011010111110",
      "001010011110001000010011001001",
      "101100001101101101100100010110",
      "011110011101001100010101111010",
      "101010011110101100000100110010",
      "000000000000010100011110110010",
      "111101100011100110000001001100",
      "100100101000101101110100000100",
      "001100111010111100101011001111",
      "000101001010101011101101010111",
      "101001011101100001100001001000",
      "001111000101101011111001000000",
      "100100010100011101100001000011",
      "000101100000101001101111000011",
      "111110010011110000100110011110",
      "011110101101011011110010110111",
      "000101100001110010001111101100",
      "111011111110111101001010010000",
      "101010110011101001111110101000",
      "001011101101001100111111111000",
      "001001011010101110110001001101",
      "101101010101001010010011100100",
      "011111011101110000010111011011",
      "011011010100001010000000011111",
      "110011001011010001010101110110",
      "100010000001010001110110000000",
      "100101111111001110011101110011",
      "110101000101000110111111111000",
      "001000100010010011110001010001",
      "001100000110101001110111010011",
      "110100101001111111110011111010",
      "001110100111111010010011011101",
      "110110110101110101001111100101",
      "110010100111011001011101100100",
      "001100100111000111100000011011",
      "101001001101001110101001100101",
      "001110101101101001110011100101",
      "100111110010011010010011000001",
      "010000101011001101110100011010",
      "101001010011111100100011100110",
      "010100011000011110111001000111",
      "000010100111110110101000001100",
      "011110000001001010000001110100",
      "000110111100000101001011101011",
      "000010010010100101000101001101",
      "101010010111101011110010010101",
      "011000101110000101011100011010",
      "001110110001111110001110000011",
      "000111011001011100011110111111",
      "001010000101001001101111110011",
      "011111000110000010100100110001",
      "011111010001101101101110011110",
      "001011011100000100101111111101",
      "100100111000011100101111110101",
      "010100011001000110010000110110",
      "011100101011010011100101001101",
      "110000111111111101011001111111",
      "001110111000101101101101101000",
      "100100110110100110011110111010",
      "011111110111100111100101101011",
      "000000001100111111110111111001",
      "101101000101111001101000100001",
      "010110000010001010001111100010",
      "100111111010111001111101110100",
      "100011110010001000011100000111",
      "000011110001011001001010111111",
      "101011111100011101010111110100",
      "111010001100111101110010101000",
      "111010000000101011110110001100",
      "011110011100110011011011101110",
      "100000111000011110001111110100",
      "001101100000100101110101011111",
      "011100101110111100011001001111",
      "110010110001001011000101001110",
      "001101101101100101000100101110",
      "011011010101100000010011101001",
      "100011101000101101100010011100",
      "001001111010100111100100100010",
      "011010100001010111111000100101",
      "000111010101101100101001110000",
      "011010100011000001001111010011",
      "110000101101101011111010001111",
      "110100100110101001101001001011",
      "101010100110001001110000101000",
      "010110100000110101011011100100",
      "000101001101100001111011110001",
      "111010001110001000001100001001",
      "000000000001110110010000110001",
      "000001000101000001000010010111",
      "011101110110101001010001110001",
      "110111000001111001010001010011",
      "011101100111110010111110010110",
      "000011000011011111011111110010",
      "001101010100100000110100110110",
      "011100111011110001001101110010",
      "010101100101110111000010000000"
    ),
    (
      "111101110100111101110111110100",
      "011111110110111100101100111111",
      "010010101011000001101110011011",
      "100010011001011001100010101001",
      "011100010000111100110111010100",
      "000110010111011101110110011010",
      "101100001101101011011000010100",
      "010110001011001110010001011001",
      "101010111101111110101010010011",
      "101100000000101011111110101001",
      "100011000100000011010110000100",
      "100001010001001101101101111111",
      "111011000001110101111111000111",
      "001001000010010010110001011001",
      "100011100010101111110001101110",
      "011001100000010001011111010000",
      "010101110001100000011111101111",
      "100000000000001000000111110010",
      "101010001111110100110010010001",
      "111101010111100110001100001110",
      "010010011111000001101101000101",
      "011001011111000011011101111010",
      "111011000000010110100110000100",
      "101011111011101101011101001010",
      "111100111110001110101101001001",
      "100101101110011100000010100001",
      "100100111010000001010010101001",
      "111110000011100101110100110000",
      "111111011011110011101100011011",
      "111100110010001011101101000110",
      "001110111011101000111110111101",
      "100010111110111010111110110000",
      "011010001001011000011101111100",
      "100110010001110001001100011001",
      "001001110100111101010011101011",
      "101011100000010001111010010111",
      "100111001000100101100001111001",
      "101110011101010110110011110001",
      "100101001110101001100010000100",
      "010000010011001111110000111010",
      "011011111011101111000010110000",
      "011100111010010110001100001100",
      "010111010111010000111011000011",
      "100111001001011100010110000011",
      "000111000010101101111101100011",
      "101001001000010110101000101101",
      "100111110001011001000010001110",
      "111110101010111010101110100101",
      "101011101110101101101001101000",
      "100001000101011010101100010111",
      "100000101101001101101001001001",
      "001000001000111110110111010100",
      "101100101100100111001011100001",
      "101010110110100001010010101000",
      "101001010000111001101100110001",
      "001101011011111111110001000010",
      "010100111000010111110101010000",
      "111010111001001010010100110000",
      "110000101001111000001111001100",
      "000100110101110111010101110001",
      "001110100010011000001100101011",
      "011000110101101001110010100011",
      "001010100100010010010010010100",
      "000101011111011100000010011010",
      "000100001010100100111011000110",
      "010001110110011101011001110001",
      "011001110111101000011010110010",
      "001101001111011000011001010110",
      "001111100100000010110001000110",
      "000111001011110010100001101010",
      "001110001011101000001000010010",
      "001010100111010010001011110001",
      "010111111011001010010001110010",
      "101001111011111110110100110011",
      "000100100011011110111100010101",
      "001100110101110011000011101101",
      "001000100100000001111001111110",
      "001001010000100011111101000110",
      "100111101110000011110100111110",
      "111100001001100101110101010101",
      "001111000010100000001101111010",
      "111011100010101101110001110111",
      "000110101001111001010100101100",
      "011001111101001000101010101011",
      "111010011000100111100011001010",
      "101010100000011010100011101110",
      "100110001111011011000011001111",
      "011001111001100110101101001011",
      "000001001100101010101000111001",
      "000001100010010111000010100111",
      "100011101011000001000010011001",
      "111001110111100110110101110010",
      "000001001010110010101000011101",
      "101110111010001111011000110101",
      "001001001011001010001101000001",
      "001100001100110001100100110100",
      "110110000010010101000101001110",
      "101100100111101101110011011011",
      "010000001001101011100001111111",
      "001110100101101111100110100111",
      "110111101011000011100100110100",
      "100110001111001000100001011010",
      "000000011101010110011000011110",
      "111010011000010111010110101111",
      "011011110000101101111100100001",
      "101100101000111110100011001111",
      "011110011101010111110100111111",
      "000110100101111101011001011011",
      "111010010011010101000011100000",
      "110000011001101001001010111101",
      "001001110010000011101001110100",
      "110001000001111100110111010100",
      "011011111000001011010110100110",
      "010100001010010111000100011001",
      "111100110111101001000111001100",
      "001111011000111000110000110100",
      "001000011001110000100000110100",
      "011011100011010100110011000011",
      "011000011110101111101010010101",
      "010001111001101000011001011000",
      "111110011100111111110101000010",
      "001010100101001101100010100111",
      "001001001101011111110110000110",
      "011010011010100100001010101001",
      "100011101011101110100111100111",
      "100101011010001000111100011111",
      "000011000100001011010001101111",
      "100010010011100011010001011110",
      "000100001111001001111101010010",
      "100000110100111001011101100001",
      "110010110100010001001101100000",
      "011110101111111000110010111101",
      "110000010001110101010110100110",
      "011010011100010000010001000110",
      "101100100101101111101001000101",
      "000010010111011100101101010001",
      "111100100111011010111111101100",
      "010111101010001111000111011101",
      "011101111111111101111101001011",
      "100111111000000000100010011100",
      "000111110111100011100000001110",
      "110001001000101111001001000011",
      "110011111000101101000000111111",
      "100000000001111000111111010101",
      "000110111010100000110010001011",
      "001101000000000110001010111011",
      "010000000100101100001110010110",
      "000010001011000000011111000111",
      "101101011101110111111010011111",
      "001110110111111000110010100100",
      "100000110000010011000010100111",
      "011011101111110111010111101001",
      "001110001001101100000011110101",
      "100001001111111010111110001001",
      "010110111001001110011111110001",
      "110110111000011101001101101110",
      "000011000110010101001111011110",
      "010000011101001000010100001100",
      "101110101010101001110111100001",
      "011100101011001011110110101010",
      "111111101111110101111110000100",
      "101000000000011100010101101011",
      "000000010100010011101100001010",
      "000111011101111110011100001010",
      "101111000101001001000100101011",
      "100001011001001110111100101111",
      "010000001101111001000010000100",
      "111011011010111100010110001001",
      "101110011100011111010111101011",
      "100000001100000001101101001110",
      "000001010010000010010010100100",
      "011011100000100011110000100111",
      "100100100011001111100000011111",
      "000011010001000000111111001011",
      "001010001101001110011111010100",
      "010101111000100100000101110010",
      "010011011000101101000010010001",
      "101111101010101100101101101000",
      "010101011110110101000101110100",
      "010000010111001001000001100001",
      "101110011001001011110000010000",
      "011110100100001011001011111111",
      "010001011101010111100101111010",
      "111011101011011100100001101110",
      "100101110100001000011000101011",
      "111100000100011001010000111001",
      "001111101100000100000001011101",
      "010101010110010011100101110110",
      "011110011100011111001011101100",
      "101101100111111111110100001001",
      "110000001101101110000011001110",
      "010101101101001101110100000100",
      "000010101001100010000101011010",
      "010001001001001111011101010010",
      "011011101001100110111011001110",
      "001010011001000000011001000101",
      "100000000100110010001001110111",
      "011110101111100001001100101010",
      "011000001101101100111100001001",
      "110101000001010110100101111101",
      "000111100101001110100000111101",
      "111111101101010100100011111101",
      "111111111001001000011000111001",
      "000110101010010100110001110000",
      "110011010100111001100100001100",
      "011001100001110100111000000001",
      "111110101101100101111110100011",
      "001101010011000000110110010110",
      "010001011101010011001111000000",
      "101000110000001010001001011100",
      "101000011000000110101101001110",
      "110111111110111100001110110001",
      "100110101101110011001001100110",
      "110010000100101100011001001001",
      "111110100011100100100111011101",
      "010001011101010111101111000110",
      "110101101110010110010001110100",
      "010100010111011001001010101010",
      "001010001010010001011110111011",
      "101110010100011100111110111011",
      "000101101010110000010001110110",
      "101110001111010111010011101000",
      "101111010011001100110101001001",
      "001110011111111010111111001111",
      "011000010001001011010001000001",
      "010100010000110000011101110000"
    ),
    (
      "000011101110001010010001000100",
      "000111000111000001001101110101",
      "001101100110110100111100101000",
      "111111011000010000101111010011",
      "111011011011110101000100001111",
      "010000101101011111101111110111",
      "001101110010110001010000110010",
      "001010100011111101110111010001",
      "101111111001110101001100101100",
      "010111001101010101110000110111",
      "011111001000100000010001001111",
      "011010101001111110100000101010",
      "110110110011001000111101111011",
      "011011111000101101000011101001",
      "101101100111010001011001011100",
      "000001111010110000100111001100",
      "101111100111100010011010010000",
      "001011111110111011011010110101",
      "011011010111011110010011100101",
      "111100100010001100111010101100",
      "101010001000101001010110000111",
      "100110010110011100110011100010",
      "010000101001111101100111000010",
      "001010100011110001110010000001",
      "010100011101111000110011110110",
      "110100111111000100000100000010",
      "101111010111110110011010001011",
      "100001110001110001100001111101",
      "011011010011001010101001010011",
      "011011011111000011010100000100",
      "000101100011010100010101100110",
      "010011111110011000011000010111",
      "000101010011101011110111001100",
      "010010111010011001110111111000",
      "110111001101100111001111101101",
      "010101101001000111001000011001",
      "111000110110010110101001000000",
      "101111111010011001000110001001",
      "100000101010100111000110011011",
      "001110100100111100101000101000",
      "010111001011111111011001100000",
      "110010110110111101001010010001",
      "101011000010100010000101111010",
      "010011101011100101101110101010",
      "001100111100011011000111100110",
      "000000111101000111100100101001",
      "000001000101010011001101011000",
      "000100110011101011001110110111",
      "000010000001010110101010111100",
      "101001111001001101110100100101",
      "101001100111011010011011011111",
      "001101000001110010111101101001",
      "111001100010000001101011001100",
      "101000100010000000011001100011",
      "111111001101101110011100000011",
      "011100001111001101100001111011",
      "110110111010000110000111011111",
      "010000111110001110000100100010",
      "101110011100110011100011010010",
      "001111011000110010100101110110",
      "110010101011111100000100010100",
      "111001001001001101001101110001",
      "100101011110010100101110011010",
      "011010100101011011111101101100",
      "111110110000111100001000101001",
      "100111110001000001010000000110",
      "011000111110110110001001010000",
      "010011010000011100001110111101",
      "010001111000101000010011001110",
      "011111101011011010111010010100",
      "110101111011111101011110111101",
      "010101000011100000010000001100",
      "011100000110011010111111001111",
      "101011001101100011100100101110",
      "111010100001001010010110100001",
      "110001010101010100001010100100",
      "001101110010010111010100111010",
      "011001001000011110110010010000",
      "100111011101000110001111111100",
      "010100010111110111111011110110",
      "011110011001010001110100001100",
      "111100101111100011110010010011",
      "100110001010011110000000000011",
      "001110111010110001111001101111",
      "111101101011000101010110101001",
      "110011010101010100001001100110",
      "101001011111011011111010011111",
      "110100001001001100110000101000",
      "111001100010101001000011110101",
      "100001100100101110111000110101",
      "010101001100001100101101100111",
      "010010010001110110101000001100",
      "100110010111001101111011010110",
      "010011010110000101000110001010",
      "000010010100110100010011001110",
      "010111001100000101000001010110",
      "011000000001100111100111110011",
      "111001101110011100010100110011",
      "001101100101100100000000101011",
      "010101111000111010011001001010",
      "101011011010001100001100110011",
      "111001011110010101010100100011",
      "100101111111110000010101110110",
      "000110010000001001000110100101",
      "011101101010011110001101110101",
      "000111001011100011000000111110",
      "000101100011011001000101101100",
      "001001000010011000001101011110",
      "000010010110000110010011011011",
      "010010100011010111000011100000",
      "011011110101110110011101011111",
      "011111000001111111011101111000",
      "110000111100011101101110111001",
      "110100110001001100101101011011",
      "101101110000100011100100101100",
      "010001010101111011010001010110",
      "101001100111111100001010110101",
      "100101110011110001000110000011",
      "011100010100011000010101101110",
      "010011111011001010010110000011",
      "101110011011100010011111010010",
      "101010110110010111000000010111",
      "110000110001110110101110101101",
      "010101111100101010110110110101",
      "010001100111011001000001011100",
      "001110011100110100100011010101",
      "110000100010010101000001110001",
      "000001000000011110000111101001",
      "000001011111110111000100110101",
      "000010110011111010110101011100",
      "010001010001011000001101101000",
      "110000001101101001110001001111",
      "000000001001101100011001011001",
      "100011100101101010100101100111",
      "110001111000011100010011111101",
      "110001110011111100011001100010",
      "011111010110011010010111110111",
      "100011001011010010010101011111",
      "000000010000001101111110010010",
      "110111001111010111111000110100",
      "000000110100100110000110111100",
      "111001100000010001111101100010",
      "111000110001101101111001000110",
      "110000000101000000111100010100",
      "101010111000100011100010010111",
      "110010111010001000001111100010",
      "001001000101100101100100011001",
      "011101100110101111110011011010",
      "000011010011111110010111011110",
      "101111011111000000011000101101",
      "000001111100011101000001100000",
      "100001001100101111110000100101",
      "101000100110100110111101110110",
      "000111010110010010111101010001",
      "011000110100100011110111001010",
      "000001100011111000100010101011",
      "011001111000100111001011111001",
      "010110010100011010110110010011",
      "010111100010111000100001111011",
      "100100010111111101101110001001",
      "010111011111000101000010101001",
      "101111001110100110001111011100",
      "101101010100011011011010001000",
      "010101000010100000010111111110",
      "111010001011100000001100101011",
      "001111101011001011111100010101",
      "001000010111111101101010100001",
      "110001101110111110110011101010",
      "000101010110010000111110000010",
      "100001011010001001000110101010",
      "011011110010100110110101001000",
      "111000110111100001000100100001",
      "101010110100001010101111111111",
      "000110000001001001101001011000",
      "110100101100100000111000101111",
      "101000111000000010000110000100",
      "011110011100100000101111101000",
      "001011001001111001001101100000",
      "101111110001111101110111101001",
      "101111000110010100100100110000",
      "001111011101001011101111001111",
      "011011000100110110011100010100",
      "101001001011001001101010111110",
      "011011011011101111000101001001",
      "111110111110011011011111000011",
      "101011110101101101100011000000",
      "001101000011110110110110101101",
      "010101100000101011101100001001",
      "110001010101010100010010111111",
      "001001100010110100100101001111",
      "111110111110010100011000010000",
      "110100010111101001101000110000",
      "010110011100110000010001000000",
      "110101111101110110001101111101",
      "111110011111001101101111101110",
      "010101000000100001100101101110",
      "011111011010001101100111110101",
      "100100111110100100101000111011",
      "100110001111001000000110011010",
      "100010001011101010000111101101",
      "101110100010100111110000110001",
      "101100110011101000000111110110",
      "100001100110000000000010101000",
      "010010010111110000001111111101",
      "010011110100110100000100000001",
      "100100101111010001001111001011",
      "000000000100110100100000001000",
      "111110111111000010001011110011",
      "011100101101011100101001001100",
      "000011001000000110101001100011",
      "001011111101100001111000010110",
      "001101000101100101010100110110",
      "010101001000110111110000011000",
      "000010011101001011101000101000",
      "110010011100011111010011001010",
      "010010000111111110111110100110",
      "000000001010111111110000110100",
      "010000001100000100100010110100",
      "001100111011011100101111010001",
      "110110101101100001101010011110",
      "100000111100000111001110110110",
      "110111101110001101101001100100",
      "001001010100000011010000110101",
      "010101100001101101110000011110",
      "101110011001101111110101100100",
      "010100001100011110000100110000"
    ),
    (
      "100111001100000111101110100010",
      "101010011100110110101000001011",
      "101101000111001011101010010100",
      "110001011110101010000101001010",
      "100111000110111110011010110001",
      "011110010010110110110000110101",
      "110010000100100101110000100011",
      "110011110001110110100001001010",
      "000010101111001110010001100100",
      "011100010110010110001011000001",
      "001110110000110000000010001001",
      "101100100101100011010101101100",
      "100101111001010101111001001110",
      "000100100000100000000100000101",
      "000101100010001101000011011010",
      "010100100011011100011001100000",
      "001100100110100010110101001110",
      "000100101101001010101001111100",
      "101101101100110110011011010000",
      "010011011110011010001100001011",
      "100011100101011001110000010110",
      "100010100000111100010010110110",
      "100110001101100000010110110011",
      "110100001110101101000000000110",
      "010111010011101000100100100100",
      "010011001000000110001101000011",
      "000101100110011101011100010010",
      "001101001101101010011001110100",
      "001111001101001111110100001101",
      "001001100101100001110001011111",
      "011101111011001000010000101110",
      "110100110000011110010101001010",
      "000111010111011100011101110001",
      "111011110010011011000001111110",
      "110011111100000100100110110010",
      "011010000010101101110111111101",
      "110101110101101110011100111101",
      "110000000011011000100000000110",
      "100100011110000000001011111101",
      "010001110000011010101111000101",
      "001001010101010100010100010100",
      "011011011100011010111011100111",
      "011001011100111100011111011011",
      "011001101011100010111110010010",
      "110011010011111111111100101011",
      "111001011101110010101000001110",
      "011001000110101000111111000111",
      "010110000111101111001101110011",
      "101110011111101010111101010110",
      "011011011111001110100101000011",
      "110111000100001101010100111000",
      "101100001101101101111010010011",
      "000001110110001110000110010011",
      "111101101100111101111000000100",
      "110100000010011100100000111000",
      "011000011010111110101000011110",
      "110011000001110000111111101000",
      "110111111111100000100101110110",
      "000111101100001010100001001010",
      "111011110010100001001001110001",
      "101000111110111011100000001000",
      "110010111101101000101010111011",
      "101011000011100100001011101110",
      "100101011000111100110011100111",
      "011001000110110110001001111101",
      "100111111101000000011010110010",
      "100111110111111011101000000101",
      "110110101111001100110010010100",
      "111010000100000010110110100000",
      "110110111000010010001000111100",
      "010101001100100101111111010100",
      "100011101101110101101111010100",
      "000001111100101101110110011010",
      "110011111100000100010100011010",
      "001011001001011101100100101011",
      "110111101100010111111001010011",
      "001111110100110110001011000010",
      "010101110001100111011100111110",
      "100010000000001110110110100011",
      "000000000110001000000110111011",
      "111110101110110010000000100111",
      "001000001100111000010001111011",
      "101101100011110110111000101110",
      "111010110000011111110110001101",
      "000000101101000010010110010000",
      "101011101100100110100111001101",
      "010011110110110011001001000011",
      "000010010100001101100010001101",
      "000100011001010010011001001010",
      "111001111011001001100000010111",
      "010010111010110110011100000010",
      "111011100010011011010001001101",
      "000001110000111001001001101001",
      "001100000110110011010100000000",
      "111001101111111101100010001001",
      "110101010100110001100110100000",
      "110111100110100010111110010001",
      "101100101101110101000111011101",
      "101011111101011010100011110000",
      "010001001100000110001110010110",
      "011011100110011011110111000110",
      "100111000100001100001001110011",
      "100011011111010010100111000101",
      "001101011101111101000011101000",
      "110100101111110111011011111111",
      "101010010111110001101111111001",
      "100001011111001110100110100111",
      "111111110111011111010111101111",
      "001000010011100001111101110110",
      "001011100001000110101010000100",
      "111111001010001001000000010101",
      "111110101110000001100011011110",
      "001100100100110110010000111101",
      "110000001101000001001110100100",
      "010111010101011111000001111001",
      "010110110100100011100110111001",
      "111011111010100110100111111100",
      "110010000111011010111001001010",
      "000010011000001110101101010011",
      "000001011010110101000011010010",
      "001101001111110110111100000111",
      "000001100101000000011011100100",
      "010101010110100010100011001010",
      "011010011111011010001100001010",
      "110100100110111000001111011001",
      "000011100000011000010101010101",
      "100010111100000100010110101011",
      "110010110111001011111111000001",
      "011100111000101110110011000001",
      "111110011011111111100011011001",
      "000110011100101111110101101100",
      "101100101001000000010111110010",
      "110010010000010001101001011000",
      "000000101111010011001010101001",
      "100101101111101101011101011101",
      "001010000001001111100100100010",
      "100101111100001100000000000011",
      "100010000110011011011101010110",
      "100001010100111011010110110011",
      "010001100011000101101011111011",
      "000111110101110010000000011000",
      "001001011111111010001010111100",
      "101110110101000010101000011001",
      "011100111100110100101001101101",
      "000000000100010110101101011111",
      "111110100110110101101010110101",
      "011100011100010101101000111110",
      "111000110100010011110111100101",
      "001010100010100000111010010000",
      "011011111001111111111100011010",
      "111000100000011000100101100101",
      "010100001001101100110111010001",
      "000100100010011011100011110101",
      "101111000000110001010011110110",
      "011101010010010111000111000001",
      "001110011100111101111000001101",
      "010000011101001011100110011111",
      "000100100100110110011110101110",
      "100100010000110110101001101100",
      "010110011001010101101101100000",
      "101000111111001101110101101011",
      "100101010101101010010101010111",
      "001001100101111110100010100000",
      "111011101101110001001101010011",
      "011110101000000010111101111000",
      "110001111100110001011010000010",
      "110000101110110100100011110001",
      "011100100101100101100100100111",
      "100010010100000000111110010111",
      "110001110110010011111110111111",
      "111010100110110001010111100010",
      "101000010001111001101110000000",
      "000110111010000110010100100110",
      "000010111001001010101010001111",
      "111001100111100111111000001101",
      "000011001011110000001110110110",
      "110010101110100001110011101111",
      "100100101010000110110011000011",
      "011001000101100101100010000001",
      "010000011100001001000001011001",
      "000011111100101101010101101110",
      "010100011000001110100011011100",
      "000001110110110011011100111001",
      "010100101101100111100100111100",
      "100011010110010010001111001110",
      "000100011001101011111111110011",
      "101010110100101011000010110101",
      "001100111010011001101000000011",
      "010000111100011001100111010101",
      "111000111110011110101101000000",
      "100111110111101110000010111101",
      "111001010111101101101100011000",
      "011001000110111011111111111100",
      "000011010100001100100111011000",
      "111000100000011000011011100100",
      "011110001100110010010101111101",
      "101010000000011010111000010100",
      "011110000111011011101011011000",
      "000011110110110101000000111110",
      "110010111101010101001010111010",
      "100101010100110011110001010000",
      "001101100101001100001011111001",
      "101110101100011010101010001101",
      "111101000000001010101111011110",
      "010101111011101000000111011011",
      "010010010101100000111001110110",
      "111010011111110101111111010110",
      "110111111000001100100111010101",
      "000011000000010000011110001010",
      "101000101000011011000111010010",
      "101111010010011001111011010001",
      "100001111101001110001001100100",
      "100001101010100000101110110011",
      "001001100000110111100110000111",
      "000001111001001100011111100001",
      "011100010001110011100011100110",
      "010101110100000110101000101100",
      "100111101100110001100001100111",
      "010011101100111010100100001100",
      "010011011100100010101010001010",
      "010010011110001010000001001101",
      "001001001010001011110111011000",
      "101010101100111101100100011010",
      "010101011100100100011110111101",
      "001011011011000111010011111001",
      "011100110111111001100100110000"
    ),
    (
      "110100111011100101100100110010",
      "100011110100110111010000100000",
      "001111111010100000101101010101",
      "100010100000010011000100110000",
      "010110110010011010001011111001",
      "010000111101010110011111101110",
      "100000000011010001111001101110",
      "100110011100100001100010111000",
      "101101111010000101100001110101",
      "010110101001111101001100100101",
      "001000100001101000001010110110",
      "001111011111001001110110001100",
      "001000010110000100101100010111",
      "100100010000100001001111110011",
      "011010100010001110101110000001",
      "111010000110000011110001001011",
      "000100111000111100100000100111",
      "011110001101011010001000100101",
      "101110100000101110101010011100",
      "111110101001111001001100110000",
      "001101100001011001110011100000",
      "110111011001111010011101100000",
      "101000100010010100110110111110",
      "101100001100111111010110111000",
      "000110111000101011010111011001",
      "010101101101110011011101011111",
      "101110101011111111111111000010",
      "010010110010010101000001101000",
      "100001110011001010101000111000",
      "000110000000001110100000100100",
      "010111111000100100110001010110",
      "000101100100010001111001011111",
      "011111000100111011000001001110",
      "101001001000110111001111001110",
      "010011100001111011011010010111",
      "010010010011010101111100110011",
      "101001100110000110100000011100",
      "100100011011110100111100100101",
      "111111000011011011110011100111",
      "100110011101100100001000100110",
      "001001101011000100101001110100",
      "100011001001100111100100001101",
      "111101111000011111001100011011",
      "001100000100100110000001011111",
      "100000000110011011011001010110",
      "001110010000001110010011010001",
      "010011000001001001111010100111",
      "010111010111000100011101110010",
      "010011110110010110111100001111",
      "110111001001010000110110010101",
      "010101010011101111101110010001",
      "101101001100000010100000101000",
      "101101100100010000010011010100",
      "101010100001110110000001001101",
      "100111110000111110101001111110",
      "001110100100001000010101010111",
      "111000000011010011101001101010",
      "000110010001101001000001010100",
      "011011011111011101001010010001",
      "111101001110001010110010010010",
      "011011100011111000101000000001",
      "111001101110000011000001001011",
      "101011001010001111000001000101",
      "000010001000011010010101011101",
      "001101110101001000001101100100",
      "010100000101110100101111001001",
      "100001101010011101000100100111",
      "110110000101111011000000111001",
      "101011010101111001000010100000",
      "001010101010000100001000011111",
      "010010011010011011000110111011",
      "111000101010001111010000111001",
      "010110111101011101001110110011",
      "101101111101000111011001010010",
      "001110000000010000010000010001",
      "101001111011011111000001011110",
      "100111111100110011011111111111",
      "101001011101101111000011100000",
      "100111100110000001011000010111",
      "111101101000010101100101000110",
      "010000110010110000100000010001",
      "111011110010100001111111100011",
      "000011101000110101010010111001",
      "010000101011000100101000110001",
      "001111000001101111000011011101",
      "100100110111100110001010110110",
      "000011000110000101000101110011",
      "001111101101001000000111101100",
      "011111111110001110111011100111",
      "011110011110100101001110001001",
      "010001010111000000000111010011",
      "111001010010100001111111111001",
      "111010010110110011100111101100",
      "111110001011110101111110100000",
      "110101110001011101010000111000",
      "111010001101000111110000010110",
      "011101011101110001110001101001",
      "000111010001000010010100111111",
      "010110101110101001000000111011",
      "110010110000000001101001001010",
      "111001100100101011001011100011",
      "100001101010111011100010111010",
      "111101101110100100101010001010",
      "100110110111111000100111001100",
      "100110111110110010011001001011",
      "001011101100000101101001011111",
      "011011010011001101000110000011",
      "001100010011111011101100110010",
      "000011111110010100011011011010",
      "110010011011000011001100011010",
      "011000101111101000010001001000",
      "100110000010100101011111001001",
      "111011100101000000110001000110",
      "101110111011001110110000110110",
      "010111010111011010100101111101",
      "100111001110000100100000110000",
      "111010001001011111101100001110",
      "000010001000101001101001110101",
      "100100111010101101110001001000",
      "110110111100111011011010100101",
      "011110001110110011011111100111",
      "011100110011101000010001011100",
      "110000001100110010010111100001",
      "111011110111111001011000110101",
      "100111101110011011110010010010",
      "101010000010001011111110000010",
      "000001111101010010000001111001",
      "010110111100010001110100100000",
      "011001011110101110111110111110",
      "010010011110111011001010100111",
      "011010101011011011001000101111",
      "100101001001111101001001100100",
      "101000010100001111000000101000",
      "010001101111000100110011011111",
      "100101010111110110101001100111",
      "011010001000011111010001101101",
      "100011000101011000100010001101",
      "101101000001101000001001011011",
      "010000000110000111101111011011",
      "000000000010000101000010100110",
      "110101100011011010011011111100",
      "100110111001101100011001011111",
      "011011011001111110110001101010",
      "011010110100101011111001100111",
      "100110011001010011111101011101",
      "011101000110110000110001101011",
      "010100100111010011001111101101",
      "111101000101101110101001100010",
      "100001111011010111001100010000",
      "101010110111110011000110101101",
      "101001101000000100110010100011",
      "001000101101100010001010010011",
      "011011100101010110100101111010",
      "011001001101100101101001101011",
      "100110101110011011101000100111",
      "011110011001101110110101001101",
      "001101110101001101100100011101",
      "000011001000010010011001101010",
      "000010010001101000001001111001",
      "110000001001010110010001111110",
      "010101110001100011011110011110",
      "111100011100100001011000010101",
      "010011010101011010011100001010",
      "001100010011001111111110110001",
      "001011111111001110010110111011",
      "101000100001011010010101110101",
      "000111110111011100111001011111",
      "111111001101001101101110010001",
      "100010100111000001001010000000",
      "001101001000001001001101010111",
      "101111101110000000011011000011",
      "000001101001011000100010001110",
      "111110011111011010110000111110",
      "011110100100101010110110011011",
      "110111000110011010000111111101",
      "000110010001101010101100001010",
      "000000001001010011010001011001",
      "110111100101100011010011100100",
      "001011111110110110000010101100",
      "010001110100101101000001100110",
      "001011110110010011010010111011",
      "011110110111101111111011110011",
      "100010100010100010101110101110",
      "001011111010110100010101010001",
      "000100000001001111110000101110",
      "011000110010110100111111000100",
      "001110010011011001100100110111",
      "111000010111111000001101010001",
      "000100010010001010001101010111",
      "010111100100010100100111001110",
      "101010010011010011000111000111",
      "101110010011011001111010000010",
      "110001001000000111001001110011",
      "111100100101110110010110101000",
      "111100001011011111110100101010",
      "001011001111000011010100010110",
      "100001010101110111010100000001",
      "010100000111111111000101001011",
      "110001000001110001100111001010",
      "000010110100010000000011101011",
      "011010011101110111010001100101",
      "101110101101000100101100111011",
      "010110111000101101111110101100",
      "000001111010010010010010111000",
      "001001110100000000111010001010",
      "000111111100110001011010000010",
      "100111110011011101110100110000",
      "110111111001100010001101011000",
      "100100011111110010111000101010",
      "001010111011110000111101110001",
      "010000001101111000110101111011",
      "001000010111111010110111100111",
      "100001100010110101110001011001",
      "001001110010000011000100001101",
      "010010001110010001000011001101",
      "010010101000001010111011100100",
      "011010111000110000001011101000",
      "111000110111100111101110000101",
      "010001001010010000101010010001",
      "000010100010101010100111010101",
      "001010110001000111110111111001",
      "110000010100001101101001010100",
      "000100110001010111010000011000",
      "000010000100100110101111000110",
      "001100010010110000101001101110",
      "000000111110110110111001100011"
    ),
    (
      "000101101011000010000001110000",
      "101101100101001001001011100000",
      "111101101011000000110011001011",
      "010100111001110110111110011010",
      "111010101110010110111110100001",
      "010111111111101111110110110010",
      "101110011111110001011000111010",
      "101001001101110111010011111110",
      "000101011100000010000001010110",
      "000011100110000111010000000010",
      "111000000000110110010000100100",
      "101110111100010000110110110110",
      "101010011101100100000001011011",
      "011011100101100010100100101101",
      "001010011101011111000010000010",
      "110101100000001001100100110110",
      "101010110001011110101011011010",
      "100001011110100001111000110101",
      "010100101011100000011101011000",
      "101011101100111011110100011110",
      "110011111001010100001111000111",
      "110101100001110010100111100000",
      "111111011001000010100000000010",
      "010100011111110110010000001100",
      "111111100101101111100010001010",
      "000001000110110000010011000010",
      "111001101110110101101100011100",
      "000111100100100100110110000100",
      "000100101011111000111011001100",
      "101011010110001011110011110110",
      "101101001000100001000001111100",
      "001110011001011001101010001010",
      "111101011100110100001111110101",
      "111011110011000001010110100110",
      "010111011111110000001110011000",
      "010100110101011100001111000010",
      "111000001110010001110101100010",
      "000000100101101001000010110000",
      "001110011010101110101110001101",
      "110011111001000101010011100110",
      "111101111100111110001000110110",
      "110001110101111001101110010011",
      "000111011011100000000000001110",
      "001000110000111011010111001101",
      "011111001101010010110100011110",
      "011010011001101110111110111011",
      "101011101001100111011001100101",
      "010101110011111001001000001111",
      "000110111000011111100101100100",
      "001001101000101001011100001001",
      "101101100111011111110100101111",
      "100011010101010101100111100100",
      "011010010110011000100011110010",
      "010000010001001010101000100111",
      "100010100111101111001011100011",
      "110100000010010100111110100011",
      "100100110001110011000000101111",
      "010001111101100111110110001110",
      "001111110101010111001101011110",
      "110000100111101001101101000111",
      "010010010101000001111111010100",
      "101010101011010001111111110111",
      "011001010110110010101100101000",
      "111000011001111110100000001010",
      "111101010111011100000101111011",
      "110101100111110100000110100111",
      "011110100000010101110110100011",
      "101111001011001111010110110101",
      "111111101100110011111011000010",
      "101100101100101101011000110001",
      "010000110111111100110011001000",
      "101000111111011011010010100001",
      "110010000001111101101110100110",
      "101010100000110111001110111110",
      "011000101011001110110011011110",
      "010001001100010011000001111001",
      "010011010111101100110111011101",
      "011011101101011000001010101001",
      "101101110111110001100010010010",
      "111001111000101111110111111110",
      "110010011001101101010010001101",
      "110101111011011101101010110110",
      "001011101010011110111010100101",
      "010000101010100000110100100011",
      "000000110010001010000001100110",
      "101000011001111111110001000110",
      "010100010111000011011111000101",
      "011001111010101001111011111011",
      "100001111010111010000000000110",
      "101111000100101110100111001010",
      "111001010110101111100111100100",
      "010110111110101100110000101111",
      "001001101100101011110110000010",
      "100100110001110010111100000100",
      "111110000010000100111111011001",
      "010010110110110110100101000100",
      "011000010000001001011111100001",
      "000110011111000001101010011011",
      "110001110100101100110010100000",
      "000101010011100100110010110111",
      "001010110000110110100110101000",
      "111100001011101101110110110010",
      "111101111100001101000100001001",
      "001111100100101100001100101111",
      "101001111001011100100100011110",
      "010101011111111100101110000111",
      "011111100000110011000011000110",
      "000001001110010000010110111000",
      "000001100000101110101001000110",
      "111011011011101101100100001011",
      "001011110111010010101011010100",
      "110100000100001111110111110000",
      "101100110000100111100001100000",
      "110001101110111101110001010100",
      "000000010111011101101000001001",
      "001101000101011100101000001010",
      "001100010001101000110101111110",
      "001100100110011011100100111010",
      "110001100011000010111110110101",
      "001010001010111100010011000001",
      "100100001010101101100001001010",
      "000010100101011010111000101100",
      "101101000010111111101010110000",
      "000100011101111010100100011010",
      "101111110100000001011000000001",
      "000010010010000111100111011100",
      "000111010000001001101100110011",
      "011001110010001101100011100010",
      "100100001101110011110001011100",
      "100000011100001010111100001000",
      "101100100001111110110011111010",
      "110010111101010010101111110010",
      "000001101111010000110111010101",
      "011000111111101001111010001110",
      "111011011100100000110011011000",
      "100000100011001110010011000000",
      "101000000101011111110010101101",
      "001001110010111101100000110100",
      "001011010000001100101101101100",
      "001111100001100001001010000110",
      "011101011111000110111001111011",
      "101010110101011010100011110010",
      "100100110110011000001010000110",
      "000100110011011100000001010101",
      "000010110011111000010100001001",
      "101010101111100100110000110001",
      "001111100010011001111010100010",
      "001001010000100000111110011000",
      "101000101001010111010011111010",
      "000010000000011101010001110111",
      "100111111111000110011110001010",
      "000111101000000110001000111101",
      "010110001110000010010111001000",
      "010101110000000110000101010101",
      "000001110001101011000010010011",
      "000101011000010110010100110010",
      "110010101101101100011011011010",
      "010010011101011101101010011100",
      "101101001110101000110101000000",
      "101001100100110101010000100011",
      "010101110100011000110101101111",
      "010110111010100100100100111110",
      "011000110100011100010111000110",
      "110101000100100000011111110111",
      "110111011011110110111010011001",
      "011100011111011000010001000011",
      "110000010000011001001100100110",
      "010001011000111001001000001000",
      "011101100100110011110101100010",
      "101101111100010000100111111011",
      "111000110000000000010110111010",
      "101100001111101101101101110001",
      "101010010111011011011000000101",
      "011000111000000100001000100100",
      "110011100010111111111100110011",
      "011111110000110000100111101011",
      "110001010101001010000110000110",
      "001011111110110110110110010101",
      "011110111101000101110010010111",
      "001100010011111110000101010110",
      "010100101011110101010110010101",
      "100101100011001111011011110010",
      "111100101100100100001100111001",
      "001110011101010110011110101111",
      "111111111000111100111101000111",
      "110010111011110010101111010001",
      "100011000011010111101101110001",
      "111000100000111011001111110111",
      "010110000010011011101001010100",
      "000010100100000001011110001010",
      "111010001001111101111000011111",
      "001010110101111101110111111100",
      "000001111110001111101110010110",
      "010001100001100000100101111000",
      "001011111001001111100100000110",
      "011111101100101001000100001000",
      "000011110110011110101010000110",
      "101000001100010111100001100000",
      "010100010000111011000100100111",
      "011110001111101110011010110100",
      "011110111101101000111011011001",
      "001101110010110010101000011111",
      "011100010010100101010101110101",
      "001111101000110100111010001111",
      "101010110101111000101000111011",
      "010100100001000110100111100010",
      "110000100011011011001000100100",
      "111111010011111100101110001100",
      "001110000101110100100100001001",
      "101001111011011000001111111010",
      "000010011100100110100110110001",
      "111101110010110100011111100001",
      "011000000101110111010011100111",
      "110111001100110100110111000101",
      "011100111100011110010001001011",
      "000110001000011011010111010101",
      "110100011111110111010101100001",
      "111000010111011011001010110000",
      "001011111111100100001100110100",
      "110010010001101000010001100001",
      "010111110100110001010100001000",
      "100110010101101110110001010100",
      "111000010111110101001100110110",
      "110000010110001011010011100101",
      "010001100011111011111111100000",
      "001011101000001110111011100000"
    )
  );

-------------------------------------------------------------------------------

  -- constants for State permutation for RMATRIX
  type INT_ARRAY is array(integer range <>) of integer;
  type R_C_ARRAY is array(0 to 5) of integer;
  type R_ARRAY is array(0 to R - 2) of R_C_ARRAY;

  -- number of columns to swap per matrix
  constant R_CC : INT_ARRAY(0 to R - 2) := (
    3,
    4,
    1,
    3,
    0,
    3,
    0,
    0,
    0,
    1,
    5,
    4,
    1,
    1,
    1,
    0,
    0,
    4,
    1,
    2,
    3,
    2,
    1,
    3,
    1,
    1,
    2,
    0,
    0,
    6,
    2,
    5,
    1,
    0,
    2,
    0,
    3
  );

  -- columns to swap per matrix
  constant R_C : R_ARRAY := (
    (
      225, 226, 227, 0, 0, 0
    ),
    (
      222, 226, 227, 228, 0, 0
    ),
    (
      223, 0, 0, 0, 0, 0
    ),
    (
      225, 226, 227, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      223, 224, 227, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      225, 0, 0, 0, 0, 0
    ),
    (
      224, 225, 226, 228, 229, 0
    ),
    (
      219, 224, 226, 228, 0, 0
    ),
    (
      224, 0, 0, 0, 0, 0
    ),
    (
      225, 0, 0, 0, 0, 0
    ),
    (
      224, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      225, 226, 227, 228, 0, 0
    ),
    (
      224, 0, 0, 0, 0, 0
    ),
    (
      224, 225, 0, 0, 0, 0
    ),
    (
      224, 226, 227, 0, 0, 0
    ),
    (
      224, 225, 0, 0, 0, 0
    ),
    (
      225, 0, 0, 0, 0, 0
    ),
    (
      221, 226, 227, 0, 0, 0
    ),
    (
      224, 0, 0, 0, 0, 0
    ),
    (
      223, 0, 0, 0, 0, 0
    ),
    (
      225, 226, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      224, 225, 226, 228, 229, 230
    ),
    (
      225, 226, 0, 0, 0, 0
    ),
    (
      222, 226, 227, 228, 229, 0
    ),
    (
      225, 0, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      225, 226, 0, 0, 0, 0
    ),
    (
      0, 0, 0, 0, 0, 0
    ),
    (
      224, 225, 226, 0, 0, 0
    )
  );

end lowmc_pkg;
